// -----------------------------------------------------------------------
//
// This is a table driven 65Cx2 core by A.Daly 
// This is a derivative of the excellent FPGA64 core see below
//
// -----------------------------------------------------------------------
// Copyright 2005-2008 by Peter Wendrich (pwsoft@syntiac.com)
// http://www.syntiac.com/fpga64.html
// -----------------------------------------------------------------------

module R65C02(
    reset,
    clk,
    enable,
    nmi_n,
    irq_n,
    di,
    dout,
    addr,
    nwe,
    sync,
    sync_irq,
    Regs
);
    
    input            reset;
    input            clk;
    input            enable;
    input            nmi_n;
    input            irq_n;
    input [7:0]      di;
    output [7:0]     dout;
    output [15:0]    addr;
    output           nwe;
    output           sync;
    output           sync_irq;
    // 6502 registers (MSB) PC, SP, P, Y, X, A (LSB)
    output [63:0]    Regs;
    
    // Store Zp    (3) => fetch, cycle2, cycleEnd
    // Store Zp,x  (4) => fetch, cycle2, preWrite, cycleEnd
    // Read  Zp,x  (4) => fetch, cycle2, cycleRead, cycleRead2
    // Rmw   Zp,x  (6) => fetch, cycle2, cycleRead, cycleRead2, cycleRmw, cycleEnd
    // Store Abs   (4) => fetch, cycle2, cycle3, cycleEnd
    // Store Abs,x (5) => fetch, cycle2, cycle3, preWrite, cycleEnd
    // Rts         (6) => fetch, cycle2, cycle3, cycleRead, cycleJump, cycleIncrEnd
    // Rti         (6) => fetch, cycle2, stack1, stack2, stack3, cycleJump
    // Jsr         (6) => fetch, cycle2, .. cycle5, cycle6, cycleJump
    // Jmp abs     (-) => fetch, cycle2, .., cycleJump
    // Jmp (ind)   (-) => fetch, cycle2, .., cycleJump
    // Brk / irq   (6) => fetch, cycle2, stack2, stack3, stack4
    // -----------------------------------------------------------------------
    
    
    //	signal counter : unsigned(27 downto 0);
    //	signal mask_irq : std_logic;
    //	signal mask_enable : std_logic;
    // Statemachine
    
    parameter [4:0]  cpuCycles_Fetch = 0,
                     cpuCycles_cycle2 = 1,
                     cpuCycles_cycle3 = 2,
                     cpuCycles_cyclePreIndirect = 3,
                     cpuCycles_cycleIndirect = 4,
                     cpuCycles_cycleBranchTaken = 5,
                     cpuCycles_cycleBranchPage = 6,
                     cpuCycles_cyclePreRead = 7,
                     cpuCycles_cycleRead = 8,
                     cpuCycles_cycleRead2 = 9,
                     cpuCycles_cycleRmw = 10,
                     cpuCycles_cyclePreWrite = 11,
                     cpuCycles_cycleWrite = 12,
                     cpuCycles_cycleStack1 = 13,
                     cpuCycles_cycleStack2 = 14,
                     cpuCycles_cycleStack3 = 15,
                     cpuCycles_cycleStack4 = 16,
                     cpuCycles_cycleJump = 17,
                     cpuCycles_cycleEnd = 18;
    // New  is read and registers updated
    // Cycle before read while doing zeropage indexed addressing.
    // Read cycle
    // Second read cycle after page-boundary crossing.
    // Calculate ALU output for read-modify-write instr.		
    // Cycle before write when doing indexed addressing.
    // Write cycle for zeropage or absolute addressing.
    // Last cycle of Jsr, Jmp. Next fetch address is target addr.
    reg [4:0]        theCpuCycle;
    reg [4:0]        nextCpuCycle;
    reg              updateRegisters;
    reg              processIrq;
    reg              nmiReg;
    reg              nmiEdge;
    reg              irqReg;		// Delay IRQ input with one clock cycle.
    wire             soReg;		// SO pin edge detection
    
    // Opcode decoding
    parameter        opcUpdateA = 0;
    parameter        opcUpdateX = 1;
    parameter        opcUpdateY = 2;
    parameter        opcUpdateS = 3;
    parameter        opcUpdateN = 4;
    parameter        opcUpdateV = 5;
    parameter        opcUpdateD = 6;
    parameter        opcUpdateI = 7;
    parameter        opcUpdateZ = 8;
    parameter        opcUpdateC = 9;
    
    parameter        opcSecondByte = 10;
    parameter        opcAbsolute = 11;
    parameter        opcZeroPage = 12;
    parameter        opcIndirect = 13;
    parameter        opcStackAddr = 14;		// Push/Pop address
    parameter        opcStackData = 15;		// Push/Pop status/data
    parameter        opcJump = 16;
    parameter        opcBranch = 17;
    parameter        indexX = 18;
    parameter        indexY = 19;
    parameter        opcStackUp = 20;
    parameter        opcWrite = 21;
    parameter        opcRmw = 22;
    parameter        opcIncrAfter = 23;		// Insert extra cycle to increment PC (RTS)
    parameter        opcRti = 24;
    parameter        opcIRQ = 25;
    
    parameter        opcInA = 26;
    parameter        opcInBrk = 27;
    parameter        opcInX = 28;
    parameter        opcInY = 29;
    parameter        opcInS = 30;
    parameter        opcInT = 31;
    parameter        opcInH = 32;
    parameter        opcInClear = 33;
    
    parameter        aluMode1From = 34;
    //
    parameter        aluMode1To = 37;
    
    parameter        aluMode2From = 38;
    //
    parameter        aluMode2To = 40;
    //
    parameter        opcInCmp = 41;
    parameter        opcInCpx = 42;
    parameter        opcInCpy = 43;
    
    //
    //               is Interrupt  -----------------+
    //          instruction is RTI ----------------+|
    //    PC++ on last cycle (RTS) ---------------+||
    //                      RMW    --------------+|||
    //                     Write   -------------+||||
    //               Pop/Stack up -------------+|||||
    //                    Branch   ---------+  ||||||
    //                      Jump ----------+|  ||||||
    //            Push or Pop data -------+||  ||||||
    //            Push or Pop addr ------+|||  ||||||
    //                   Indirect  -----+||||  ||||||
    //                    ZeroPage ----+|||||  ||||||
    //                    Absolute ---+||||||  ||||||
    //              PC++ on cycle2 --+|||||||  ||||||
    //                               |AZI||JBXY|WM|||
    parameter [0:15] immediate = 16'b1000000000000000;
    parameter [0:15] implied = 16'b0000000000000000;
    // Zero page
    parameter [0:15] readZp = 16'b1010000000000000;
    parameter [0:15] writeZp = 16'b1010000000010000;
    parameter [0:15] rmwZp = 16'b1010000000001000;
    // Zero page indexed
    parameter [0:15] readZpX = 16'b1010000010000000;
    parameter [0:15] writeZpX = 16'b1010000010010000;
    parameter [0:15] rmwZpX = 16'b1010000010001000;
    parameter [0:15] readZpY = 16'b1010000001000000;
    parameter [0:15] writeZpY = 16'b1010000001010000;
    parameter [0:15] rmwZpY = 16'b1010000001001000;
    // Zero page indirect
    parameter [0:15] readIndX = 16'b1001000010000000;
    parameter [0:15] writeIndX = 16'b1001000010010000;
    parameter [0:15] rmwIndX = 16'b1001000010001000;
    parameter [0:15] readIndY = 16'b1001000001000000;
    parameter [0:15] writeIndY = 16'b1001000001010000;
    parameter [0:15] rmwIndY = 16'b1001000001001000;
    parameter [0:15] rmwInd = 16'b1001000000001000;
    parameter [0:15] readInd = 16'b1001000000000000;
    parameter [0:15] writeInd = 16'b1001000000010000;
    //                               |AZI||JBXY|WM||
    // Absolute
    parameter [0:15] readAbs = 16'b1100000000000000;
    parameter [0:15] writeAbs = 16'b1100000000010000;
    parameter [0:15] rmwAbs = 16'b1100000000001000;
    parameter [0:15] readAbsX = 16'b1100000010000000;
    parameter [0:15] writeAbsX = 16'b1100000010010000;
    parameter [0:15] rmwAbsX = 16'b1100000010001000;
    parameter [0:15] readAbsY = 16'b1100000001000000;
    parameter [0:15] writeAbsY = 16'b1100000001010000;
    parameter [0:15] rmwAbsY = 16'b1100000001001000;
    // PHA PHP
    parameter [0:15] push = 16'b0000010000000000;
    // PLA PLP
    parameter [0:15] pop = 16'b0000010000100000;
    // Jumps
    parameter [0:15] jsr = 16'b1000101000000000;
    parameter [0:15] jumpAbs = 16'b1000001000000000;
    parameter [0:15] jumpInd = 16'b1100001000000000;
    parameter [0:15] jumpIndX = 16'b1100001010000000;
    parameter [0:15] relative = 16'b1000000100000000;
    // Specials
    parameter [0:15] rts = 16'b0000101000100100;
    parameter [0:15] rti = 16'b0000111000100010;
    parameter [0:15] brk = 16'b1000111000000001;
    //	constant irq       : addrDef $ "0000111000000001";
    //	constant        : unsigned(0 to 0) $ "0";
    parameter [0:15] xxxxxxxx = 16'bxxxxxxxxxx0xxx00;
    
    // A = accu
    // X = index X
    // Y = index Y
    // S = Stack pointer
    // H = indexH
    // 
    //                                       AEXYSTHc
    parameter [0:7]  aluInA = 8'b10000000;
    parameter [0:7]  aluInBrk = 8'b01000000;
    parameter [0:7]  aluInX = 8'b00100000;
    parameter [0:7]  aluInY = 8'b00010000;
    parameter [0:7]  aluInS = 8'b00001000;
    parameter [0:7]  aluInT = 8'b00000100;
    parameter [0:7]  aluInClr = 8'b00000001;
    parameter [0:7]  aluInSet = 8'b00000000;
    parameter [0:7]  aluInXXX = 8'bxxxxxxxx;
    
    // Most of the aluModes are just like the s.
    // aluModeInp -> input is output. calculate N and Z
    // aluModeCmp -> Compare for CMP, CPX, CPY
    // aluModeFlg -> input to flags needed for PLP, RTI and CLC, SEC, CLV
    // aluModeInc -> for INC but also INX, INY
    // aluModeDec -> for DEC but also DEX, DEY
    
    
    // Logic/Shift ALU
    parameter [0:3]  aluModeInp = 4'b0000;
    parameter [0:3]  aluModeP = 4'b0001;
    parameter [0:3]  aluModeInc = 4'b0010;
    parameter [0:3]  aluModeDec = 4'b0011;
    parameter [0:3]  aluModeFlg = 4'b0100;
    parameter [0:3]  aluModeBit = 4'b0101;
    // 0110
    // 0111
    parameter [0:3]  aluModeLsr = 4'b1000;
    parameter [0:3]  aluModeRor = 4'b1001;
    parameter [0:3]  aluModeAsl = 4'b1010;
    parameter [0:3]  aluModeRol = 4'b1011;
    parameter [0:3]  aluModeTSB = 4'b1100;
    parameter [0:3]  aluModeTRB = 4'b1101;
    // 1110
    // 1111;
    
    // Arithmetic ALU
    parameter [0:2]  aluModePss = 3'b000;
    parameter [0:2]  aluModeCmp = 3'b001;
    parameter [0:2]  aluModeAdc = 3'b010;
    parameter [0:2]  aluModeSbc = 3'b011;
    parameter [0:2]  aluModeAnd = 3'b100;
    parameter [0:2]  aluModeOra = 3'b101;
    parameter [0:2]  aluModeEor = 3'b110;
    parameter [0:2]  aluModeNoF = 3'b111;
    //aluModeBRK
    //constant aluBrk  : aluMode $ aluModeBRK & aluModePss & "---";
    //constant aluFix  : aluMode $ aluModeInp & aluModeNoF & "---";
    parameter [0:9]  aluInp = {aluModeInp, aluModePss, 3'bxxx};
    parameter [0:9]  aluP = {aluModeP, aluModePss, 3'bxxx};
    parameter [0:9]  aluInc = {aluModeInc, aluModePss, 3'bxxx};
    parameter [0:9]  aluDec = {aluModeDec, aluModePss, 3'bxxx};
    parameter [0:9]  aluFlg = {aluModeFlg, aluModePss, 3'bxxx};
    parameter [0:9]  aluBit = {aluModeBit, aluModeAnd, 3'bxxx};
    parameter [0:9]  aluRor = {aluModeRor, aluModePss, 3'bxxx};
    parameter [0:9]  aluLsr = {aluModeLsr, aluModePss, 3'bxxx};
    parameter [0:9]  aluRol = {aluModeRol, aluModePss, 3'bxxx};
    parameter [0:9]  aluAsl = {aluModeAsl, aluModePss, 3'bxxx};
    parameter [0:9]  aluTSB = {aluModeTSB, aluModePss, 3'bxxx};
    parameter [0:9]  aluTRB = {aluModeTRB, aluModePss, 3'bxxx};
    parameter [0:9]  aluCmp = {aluModeInp, aluModeCmp, 3'b100};
    parameter [0:9]  aluCpx = {aluModeInp, aluModeCmp, 3'b010};
    parameter [0:9]  aluCpy = {aluModeInp, aluModeCmp, 3'b001};
    parameter [0:9]  aluAdc = {aluModeInp, aluModeAdc, 3'bxxx};
    parameter [0:9]  aluSbc = {aluModeInp, aluModeSbc, 3'bxxx};
    parameter [0:9]  aluAnd = {aluModeInp, aluModeAnd, 3'bxxx};
    parameter [0:9]  aluOra = {aluModeInp, aluModeOra, 3'bxxx};
    parameter [0:9]  aluEor = {aluModeInp, aluModeEor, 3'bxxx};
    
    parameter [0:9]  aluXXX = 1'bx;
    
    // Stack operations. Push/Pop/None
    parameter [0:0]  stackInc = 1'b0;
    parameter [0:0]  stackDec = 1'b1;
    parameter [0:0]  stackXXX = 1'bx;
    
    // +------- Update register A
    // |+------ Update register X
    // ||+----- Update register Y
    // |||+---- Update register S
    // ||||       +-- Update Flags
    // ||||       |   
    // ||||      _|__ 
    // ||||     /    \
    // AXYS     NVDIZC    addressing  aluInput  aluMode
    // AXYS     NVDIZC    addressing  aluInput  aluMode  
    // 00 BRK
    // 01 ORA (zp,x)
    // 02 NOP ------- 65C02
    // 03 NOP ------- 65C02
    // 04 TSB zp ----------- 65C02
    // 05 ORA zp
    // 06 ASL zp
    // 07 NOP ------- 65C02
    // 08 PHP
    // 09 ORA imm
    // 0A ASL accu
    // 0B NOP ------- 65C02
    // 0C TSB abs ---------- 65C02
    // 0D ORA abs
    // 0E ASL abs
    // 0F NOP ------- 65C02
    // 10 BPL
    // 11 ORA (zp),y
    // 12 ORA (zp) --------- 65C02  
    // 13 NOP ------- 65C02
    // 14 TRB zp ~---------- 65C02 
    // 15 ORA zp,x
    // 16 ASL zp,x
    // 17 NOP ------- 65C02
    // 18 CLC
    // 19 ORA abs,y
    // 1A INC accu --------- 65C02
    // 1B NOP ------- 65C02
    // 1C TRB abs ~----- --- 65C02 
    // 1D ORA abs,x
    // 1E ASL abs,x
    // 1F NOP ------- 65C02
    // AXYS     NVDIZC    addressing  aluInput  aluMode
    // 20 JSR
    // 21 AND (zp,x)
    // 22 NOP ------- 65C02
    // 23 NOP ------- 65C02
    // 24 BIT zp
    // 25 AND zp
    // 26 ROL zp
    // 27 NOP ------- 65C02
    // 28 PLP
    // 29 AND imm
    // 2A ROL accu
    // 2B NOP ------- 65C02
    // 2C BIT abs
    // 2D AND abs
    // 2E ROL abs
    // 2F NOP ------- 65C02
    // 30 BMI
    // 31 AND (zp),y
    // 32 AND (zp) -------- 65C02 
    // 33 NOP ------- 65C02
    // 34 BIT zp,x -------- 65C02
    // 35 AND zp,x
    // 36 ROL zp,x
    // 37 NOP ------- 65C02
    // 38 SEC
    // 39 AND abs,y
    // 3A DEC accu -------- 65C12
    // 3B NOP ------- 65C02
    // 3C BIT abs,x ------- 65C02
    // 3D AND abs,x
    // 3E ROL abs,x
    // 3F NOP ------- 65C02
    // AXYS     NVDIZC    addressing  aluInput  aluMode
    // 40 RTI
    // 41 EOR (zp,x)
    // 42 NOP ------- 65C02
    // 43 NOP ------- 65C02
    // 44 NOP ------- 65C02
    // 45 EOR zp
    // 46 LSR zp
    // 47 NOP ------- 65C02
    // 48 PHA
    // 49 EOR imm
    // 4A LSR accu -------- 65C02
    // 4B NOP ------- 65C02
    // 4C JMP abs
    // 4D EOR abs
    // 4E LSR abs
    // 4F NOP ------- 65C02
    // 50 BVC
    // 51 EOR (zp),y
    // 52 EOR (zp) -------- 65C02 
    // 53 NOP ------- 65C02
    // 54 NOP ------- 65C02
    // 55 EOR zp,x
    // 56 LSR zp,x
    // 57 NOP ------- 65C02
    // 58 CLI
    // 59 EOR abs,y
    // 5A PHY ------------- 65C02
    // 5B NOP ------- 65C02
    // 5C NOP ------- 65C02
    // 5D EOR abs,x
    // 5E LSR abs,x
    // 5F NOP ------- 65C02
    // AXYS     NVDIZC    addressing  aluInput  aluMode
    // 60 RTS
    // 61 ADC (zp,x)
    // 62 NOP ------- 65C02
    // 63 NOP ------- 65C02
    // 64 STZ zp ---------- 65C02
    // 65 ADC zp
    // 66 ROR zp
    // 67 NOP ------- 65C02
    // 68 PLA
    // 69 ADC imm
    // 6A ROR accu
    // 6B NOP ------ 65C02
    // 6C JMP indirect
    // 6D ADC abs
    // 6E ROR abs
    // 6F NOP ------ 65C02
    // 70 BVS
    // 71 ADC (zp),y
    // 72 ADC (zp) -------- 65C02 
    // 73 NOP ------ 65C02
    // 74 STZ zp,x -------- 65C02
    // 75 ADC zp,x
    // 76 ROR zp,x
    // 77 NOP ----- 65C02
    // 78 SEI
    // 79 ADC abs,y
    // 7A PLY ------------- 65C02
    // 7B NOP ----- 65C02
    // 7C JMP indirect,x -- 65C02
    //"0000" & "000000" & jumpInd   & aluInXXX & aluXXX, -- 6C JMP indirect
    // 7D ADC abs,x
    // 7E ROR abs,x
    // 7F NOP ----- 65C02
    // AXYS     NVDIZC    addressing  aluInput  aluMode
    // 80 BRA ----------- 65C02
    // 81 STA (zp,x)
    // 82 NOP ----- 65C02
    // 83 NOP ----- 65C02
    // 84 STY zp
    // 85 STA zp
    // 86 STX zp
    // 87 NOP ----- 65C02
    // 88 DEY
    // 89 BIT imm ------- 65C02
    // 8A TXA
    // 8B NOP ----- 65C02
    // 8C STY abs ------- 65C02
    // 8D STA abs
    // 8E STX abs
    // 8F NOP ----- 65C02
    // 90 BCC
    // 91 STA (zp),y
    // 92 STA (zp) ------ 65C02 
    // 93 NOP ----- 65C02
    // 94 STY zp,x
    // 95 STA zp,x
    // 96 STX zp,y
    // 97 NOP ----- 65C02
    // 98 TYA
    // 99 STA abs,y
    // 9A TXS
    // 9B NOP ----- 65C02
    // 9C STZ Abs ------- 65C02
    // 9D STA abs,x
    // 9C STZ Abs,x ----- 65C02
    // 9F NOP ----- 65C02
    // AXYS     NVDIZC    addressing  aluInput  aluMode
    // A0 LDY imm
    // A1 LDA (zp,x)
    // A2 LDX imm
    // A3 NOP ----- 65C02
    // A4 LDY zp
    // A5 LDA zp
    // A6 LDX zp
    // A7 NOP ----- 65C02
    // A8 TAY
    // A9 LDA imm
    // AA TAX
    // AB NOP ----- 65C02
    // AC LDY abs
    // AD LDA abs
    // AE LDX abs
    // AF NOP ----- 65C02
    // B0 BCS
    // B1 LDA (zp),y
    // B2 LDA (zp) ------ 65C02 
    // B3 NOP ----- 65C02
    // B4 LDY zp,x
    // B5 LDA zp,x
    // B6 LDX zp,y
    // B7 NOP ----- 65C02
    // B8 CLV
    // B9 LDA abs,y
    // BA TSX
    // BB NOP ----- 65C02
    // BC LDY abs,x
    // BD LDA abs,x
    // BE LDX abs,y
    // BF NOP ----- 65C02
    // AXYS     NVDIZC    addressing  aluInput  aluMode
    // C0 CPY imm
    // C1 CMP (zp,x)
    // C2 NOP ----- 65C02
    // C3 NOP ----- 65C02
    // C4 CPY zp
    // C5 CMP zp
    // C6 DEC zp
    // C7 NOP ----- 65C02
    // C8 INY
    // C9 CMP imm
    // CA DEX
    // CB NOP ----- 65C02
    // CC CPY abs
    // CD CMP abs
    // CE DEC abs
    // CF NOP ----- 65C02
    // D0 BNE
    // D1 CMP (zp),y
    // D2 CMP (zp) ------ 65C02 
    // D3 NOP ----- 65C02
    // D4 NOP ----- 65C02
    // D5 CMP zp,x
    // D6 DEC zp,x
    // D7 NOP ----- 65C02
    // D8 CLD
    // D9 CMP abs,y
    // DA PHX ----------- 65C02
    // DB NOP ----- 65C02
    // DC NOP ----- 65C02
    // DD CMP abs,x
    // DE DEC abs,x
    // DF NOP ----- 65C02
    // AXYS    NVDIZC    addressing  aluInput  aluMode
    // E0 CPX imm
    // E1 SBC (zp,x)
    // E2 NOP ----- 65C02
    // E3 NOP ----- 65C02
    // E4 CPX zp
    // E5 SBC zp
    // E6 INC zp
    // E7 NOP ----- 65C02
    // E8 INX
    // E9 SBC imm
    // EA NOP
    // EB NOP ----- 65C02
    // EC CPX abs
    // ED SBC abs
    // EE INC abs
    // EF NOP ----- 65C02
    // F0 BEQ
    // F1 SBC (zp),y
    // F2 SBC (zp) ------ 65C02 
    // F3 NOP ----- 65C02
    // F4 NOP ----- 65C02
    // F5 SBC zp,x
    // F6 INC zp,x
    // F7 NOP  ---- 65C02
    // F8 SED
    // F9 SBC abs,y
    // FA PLX ----------- 65C02
    // FB NOP ----- 65C02
    // FC NOP ----- 65C02
    // FD SBC abs,x
    // FE INC abs,x
   
    
    reg [0:43] InfoTable[255];
    initial
    begin

InfoTable[0] = {4'b0000, 6'b001100, brk, aluInBrk, aluP};
InfoTable[1] = {4'b1000, 6'b100010, readIndX, aluInT, aluOra};
InfoTable[2] = {4'b0000, 6'b000000, immediate, aluInXXX, aluXXX};
InfoTable[3] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[4] = {4'b0000, 6'b000010, rmwZp, aluInT, aluTSB};
InfoTable[5] = {4'b1000, 6'b100010, readZp, aluInT, aluOra};
InfoTable[6] = {4'b0000, 6'b100011, rmwZp, aluInT, aluAsl};
InfoTable[7] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[8] = {4'b0000, 6'b000000, push, aluInXXX, aluP};
InfoTable[9] = {4'b1000, 6'b100010, immediate, aluInT, aluOra};
InfoTable[10] = {4'b1000, 6'b100011, implied, aluInA, aluAsl};
InfoTable[11] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[12] = {4'b0000, 6'b000010, rmwAbs, aluInT, aluTSB};
InfoTable[13] = {4'b1000, 6'b100010, readAbs, aluInT, aluOra};
InfoTable[14] = {4'b0000, 6'b100011, rmwAbs, aluInT, aluAsl};
InfoTable[15] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[16] = {4'b0000, 6'b000000, relative, aluInXXX, aluXXX};
InfoTable[17] = {4'b1000, 6'b100010, readIndY, aluInT, aluOra};
InfoTable[18] = {4'b1000, 6'b100010, readInd, aluInT, aluOra};
InfoTable[19] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[20] = {4'b0000, 6'b000010, rmwZp, aluInT, aluTRB};
InfoTable[21] = {4'b1000, 6'b100010, readZpX, aluInT, aluOra};
InfoTable[22] = {4'b0000, 6'b100011, rmwZpX, aluInT, aluAsl};
InfoTable[23] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[24] = {4'b0000, 6'b000001, implied, aluInClr, aluFlg};
InfoTable[25] = {4'b1000, 6'b100010, readAbsY, aluInT, aluOra};
InfoTable[26] = {4'b1000, 6'b100010, implied, aluInA, aluInc};
InfoTable[27] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[28] = {4'b0000, 6'b000010, rmwAbs, aluInT, aluTRB};
InfoTable[29] = {4'b1000, 6'b100010, readAbsX, aluInT, aluOra};
InfoTable[30] = {4'b0000, 6'b100011, rmwAbsX, aluInT, aluAsl};
InfoTable[31] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[32] = {4'b0000, 6'b000000, jsr, aluInXXX, aluXXX};
InfoTable[33] = {4'b1000, 6'b100010, readIndX, aluInT, aluAnd};
InfoTable[34] = {4'b0000, 6'b000000, immediate, aluInXXX, aluXXX};
InfoTable[35] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[36] = {4'b0000, 6'b110010, readZp, aluInT, aluBit};
InfoTable[37] = {4'b1000, 6'b100010, readZp, aluInT, aluAnd};
InfoTable[38] = {4'b0000, 6'b100011, rmwZp, aluInT, aluRol};
InfoTable[39] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[40] = {4'b0000, 6'b111111, pop, aluInT, aluFlg};
InfoTable[41] = {4'b1000, 6'b100010, immediate, aluInT, aluAnd};
InfoTable[42] = {4'b1000, 6'b100011, implied, aluInA, aluRol};
InfoTable[43] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[44] = {4'b0000, 6'b110010, readAbs, aluInT, aluBit};
InfoTable[45] = {4'b1000, 6'b100010, readAbs, aluInT, aluAnd};
InfoTable[46] = {4'b0000, 6'b100011, rmwAbs, aluInT, aluRol};
InfoTable[47] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[48] = {4'b0000, 6'b000000, relative, aluInXXX, aluXXX};
InfoTable[49] = {4'b1000, 6'b100010, readIndY, aluInT, aluAnd};
InfoTable[50] = {4'b1000, 6'b100010, readInd, aluInT, aluAnd};
InfoTable[51] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[52] = {4'b0000, 6'b110010, readZpX, aluInT, aluBit};
InfoTable[53] = {4'b1000, 6'b100010, readZpX, aluInT, aluAnd};
InfoTable[54] = {4'b0000, 6'b100011, rmwZpX, aluInT, aluRol};
InfoTable[55] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[56] = {4'b0000, 6'b000001, implied, aluInSet, aluFlg};
InfoTable[57] = {4'b1000, 6'b100010, readAbsY, aluInT, aluAnd};
InfoTable[58] = {4'b1000, 6'b100010, implied, aluInA, aluDec};
InfoTable[59] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[60] = {4'b0000, 6'b110010, readAbsX, aluInT, aluBit};
InfoTable[61] = {4'b1000, 6'b100010, readAbsX, aluInT, aluAnd};
InfoTable[62] = {4'b0000, 6'b100011, rmwAbsX, aluInT, aluRol};
InfoTable[63] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[64] = {4'b0000, 6'b111111, rti, aluInT, aluFlg};
InfoTable[65] = {4'b1000, 6'b100010, readIndX, aluInT, aluEor};
InfoTable[66] = {4'b0000, 6'b000000, immediate, aluInXXX, aluXXX};
InfoTable[67] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[68] = {4'b0000, 6'b000000, immediate, aluInXXX, aluXXX};
InfoTable[69] = {4'b1000, 6'b100010, readZp, aluInT, aluEor};
InfoTable[70] = {4'b0000, 6'b100011, rmwZp, aluInT, aluLsr};
InfoTable[71] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[72] = {4'b0000, 6'b000000, push, aluInA, aluInp};
InfoTable[73] = {4'b1000, 6'b100010, immediate, aluInT, aluEor};
InfoTable[74] = {4'b1000, 6'b100011, implied, aluInA, aluLsr};
InfoTable[75] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[76] = {4'b0000, 6'b000000, jumpAbs, aluInXXX, aluXXX};
InfoTable[77] = {4'b1000, 6'b100010, readAbs, aluInT, aluEor};
InfoTable[78] = {4'b0000, 6'b100011, rmwAbs, aluInT, aluLsr};
InfoTable[79] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[80] = {4'b0000, 6'b000000, relative, aluInXXX, aluXXX};
InfoTable[81] = {4'b1000, 6'b100010, readIndY, aluInT, aluEor};
InfoTable[82] = {4'b1000, 6'b100010, readInd, aluInT, aluEor};
InfoTable[83] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[84] = {4'b0000, 6'b000000, immediate, aluInXXX, aluXXX};
InfoTable[85] = {4'b1000, 6'b100010, readZpX, aluInT, aluEor};
InfoTable[86] = {4'b0000, 6'b100011, rmwZpX, aluInT, aluLsr};
InfoTable[87] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[88] = {4'b0000, 6'b000100, implied, aluInClr, aluXXX};
InfoTable[89] = {4'b1000, 6'b100010, readAbsY, aluInT, aluEor};
InfoTable[90] = {4'b0000, 6'b000000, push, aluInY, aluInp};
InfoTable[91] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[92] = {4'b0000, 6'b000000, readAbs, aluInXXX, aluXXX};
InfoTable[93] = {4'b1000, 6'b100010, readAbsX, aluInT, aluEor};
InfoTable[94] = {4'b0000, 6'b100011, rmwAbsX, aluInT, aluLsr};
InfoTable[95] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[96] = {4'b0000, 6'b000000, rts, aluInXXX, aluXXX};
InfoTable[97] = {4'b1000, 6'b110011, readIndX, aluInT, aluAdc};
InfoTable[98] = {4'b0000, 6'b000000, immediate, aluInXXX, aluXXX};
InfoTable[99] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[100] = {4'b0000, 6'b000000, writeZp, aluInClr, aluInp};
InfoTable[101] = {4'b1000, 6'b110011, readZp, aluInT, aluAdc};
InfoTable[102] = {4'b0000, 6'b100011, rmwZp, aluInT, aluRor};
InfoTable[103] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[104] = {4'b1000, 6'b100010, pop, aluInT, aluInp};
InfoTable[105] = {4'b1000, 6'b110011, immediate, aluInT, aluAdc};
InfoTable[106] = {4'b1000, 6'b100011, implied, aluInA, aluRor};
InfoTable[107] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[108] = {4'b0000, 6'b000000, jumpInd, aluInXXX, aluXXX};
InfoTable[109] = {4'b1000, 6'b110011, readAbs, aluInT, aluAdc};
InfoTable[110] = {4'b0000, 6'b100011, rmwAbs, aluInT, aluRor};
InfoTable[111] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[112] = {4'b0000, 6'b000000, relative, aluInXXX, aluXXX};
InfoTable[113] = {4'b1000, 6'b110011, readIndY, aluInT, aluAdc};
InfoTable[114] = {4'b1000, 6'b110011, readInd, aluInT, aluAdc};
InfoTable[115] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[116] = {4'b0000, 6'b000000, writeZpX, aluInClr, aluInp};
InfoTable[117] = {4'b1000, 6'b110011, readZpX, aluInT, aluAdc};
InfoTable[118] = {4'b0000, 6'b100011, rmwZpX, aluInT, aluRor};
InfoTable[119] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[120] = {4'b0000, 6'b000100, implied, aluInSet, aluXXX};
InfoTable[121] = {4'b1000, 6'b110011, readAbsY, aluInT, aluAdc};
InfoTable[122] = {4'b0010, 6'b100010, pop, aluInT, aluInp};
InfoTable[123] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[124] = {4'b0000, 6'b000000, jumpIndX, aluInXXX, aluXXX};
InfoTable[125] = {4'b1000, 6'b110011, readAbsX, aluInT, aluAdc};
InfoTable[126] = {4'b0000, 6'b100011, rmwAbsX, aluInT, aluRor};
InfoTable[127] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[128] = {4'b0000, 6'b000000, relative, aluInXXX, aluXXX};
InfoTable[129] = {4'b0000, 6'b000000, writeIndX, aluInA, aluInp};
InfoTable[130] = {4'b0000, 6'b000000, immediate, aluInXXX, aluXXX};
InfoTable[131] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[132] = {4'b0000, 6'b000000, writeZp, aluInY, aluInp};
InfoTable[133] = {4'b0000, 6'b000000, writeZp, aluInA, aluInp};
InfoTable[134] = {4'b0000, 6'b000000, writeZp, aluInX, aluInp};
InfoTable[135] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[136] = {4'b0010, 6'b100010, implied, aluInY, aluDec};
InfoTable[137] = {4'b0000, 6'b000010, immediate, aluInT, aluBit};
InfoTable[138] = {4'b1000, 6'b100010, implied, aluInX, aluInp};
InfoTable[139] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[140] = {4'b0000, 6'b000000, writeAbs, aluInY, aluInp};
InfoTable[141] = {4'b0000, 6'b000000, writeAbs, aluInA, aluInp};
InfoTable[142] = {4'b0000, 6'b000000, writeAbs, aluInX, aluInp};
InfoTable[143] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[144] = {4'b0000, 6'b000000, relative, aluInXXX, aluXXX};
InfoTable[145] = {4'b0000, 6'b000000, writeIndY, aluInA, aluInp};
InfoTable[146] = {4'b0000, 6'b000000, writeInd, aluInA, aluInp};
InfoTable[147] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[148] = {4'b0000, 6'b000000, writeZpX, aluInY, aluInp};
InfoTable[149] = {4'b0000, 6'b000000, writeZpX, aluInA, aluInp};
InfoTable[150] = {4'b0000, 6'b000000, writeZpY, aluInX, aluInp};
InfoTable[151] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[152] = {4'b1000, 6'b100010, implied, aluInY, aluInp};
InfoTable[153] = {4'b0000, 6'b000000, writeAbsY, aluInA, aluInp};
InfoTable[154] = {4'b0001, 6'b000000, implied, aluInX, aluInp};
InfoTable[155] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[156] = {4'b0000, 6'b000000, writeAbs, aluInClr, aluInp};
InfoTable[157] = {4'b0000, 6'b000000, writeAbsX, aluInA, aluInp};
InfoTable[158] = {4'b0000, 6'b000000, writeAbsX, aluInClr, aluInp};
InfoTable[159] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[160] = {4'b0010, 6'b100010, immediate, aluInT, aluInp};
InfoTable[161] = {4'b1000, 6'b100010, readIndX, aluInT, aluInp};
InfoTable[162] = {4'b0100, 6'b100010, immediate, aluInT, aluInp};
InfoTable[163] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[164] = {4'b0010, 6'b100010, readZp, aluInT, aluInp};
InfoTable[165] = {4'b1000, 6'b100010, readZp, aluInT, aluInp};
InfoTable[166] = {4'b0100, 6'b100010, readZp, aluInT, aluInp};
InfoTable[167] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[168] = {4'b0010, 6'b100010, implied, aluInA, aluInp};
InfoTable[169] = {4'b1000, 6'b100010, immediate, aluInT, aluInp};
InfoTable[170] = {4'b0100, 6'b100010, implied, aluInA, aluInp};
InfoTable[171] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[172] = {4'b0010, 6'b100010, readAbs, aluInT, aluInp};
InfoTable[173] = {4'b1000, 6'b100010, readAbs, aluInT, aluInp};
InfoTable[174] = {4'b0100, 6'b100010, readAbs, aluInT, aluInp};
InfoTable[175] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[176] = {4'b0000, 6'b000000, relative, aluInXXX, aluXXX};
InfoTable[177] = {4'b1000, 6'b100010, readIndY, aluInT, aluInp};
InfoTable[178] = {4'b1000, 6'b100010, readInd, aluInT, aluInp};
InfoTable[179] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[180] = {4'b0010, 6'b100010, readZpX, aluInT, aluInp};
InfoTable[181] = {4'b1000, 6'b100010, readZpX, aluInT, aluInp};
InfoTable[182] = {4'b0100, 6'b100010, readZpY, aluInT, aluInp};
InfoTable[183] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[184] = {4'b0000, 6'b010000, implied, aluInClr, aluFlg};
InfoTable[185] = {4'b1000, 6'b100010, readAbsY, aluInT, aluInp};
InfoTable[186] = {4'b0100, 6'b100010, implied, aluInS, aluInp};
InfoTable[187] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[188] = {4'b0010, 6'b100010, readAbsX, aluInT, aluInp};
InfoTable[189] = {4'b1000, 6'b100010, readAbsX, aluInT, aluInp};
InfoTable[190] = {4'b0100, 6'b100010, readAbsY, aluInT, aluInp};
InfoTable[191] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[192] = {4'b0000, 6'b100011, immediate, aluInT, aluCpy};
InfoTable[193] = {4'b0000, 6'b100011, readIndX, aluInT, aluCmp};
InfoTable[194] = {4'b0000, 6'b000000, immediate, aluInXXX, aluXXX};
InfoTable[195] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[196] = {4'b0000, 6'b100011, readZp, aluInT, aluCpy};
InfoTable[197] = {4'b0000, 6'b100011, readZp, aluInT, aluCmp};
InfoTable[198] = {4'b0000, 6'b100010, rmwZp, aluInT, aluDec};
InfoTable[199] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[200] = {4'b0010, 6'b100010, implied, aluInY, aluInc};
InfoTable[201] = {4'b0000, 6'b100011, immediate, aluInT, aluCmp};
InfoTable[202] = {4'b0100, 6'b100010, implied, aluInX, aluDec};
InfoTable[203] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[204] = {4'b0000, 6'b100011, readAbs, aluInT, aluCpy};
InfoTable[204] = {4'b0000, 6'b100011, readAbs, aluInT, aluCmp};
InfoTable[205] = {4'b0000, 6'b100010, rmwAbs, aluInT, aluDec};
InfoTable[206] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[207] = {4'b0000, 6'b000000, relative, aluInXXX, aluXXX};
InfoTable[208] = {4'b0000, 6'b100011, readIndY, aluInT, aluCmp};
InfoTable[209] = {4'b0000, 6'b100011, readInd, aluInT, aluCmp};
InfoTable[210] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[211] = {4'b0000, 6'b000000, immediate, aluInXXX, aluXXX};
InfoTable[212] = {4'b0000, 6'b100011, readZpX, aluInT, aluCmp};
InfoTable[213] = {4'b0000, 6'b100010, rmwZpX, aluInT, aluDec};
InfoTable[214] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[215] = {4'b0000, 6'b001000, implied, aluInClr, aluXXX};
InfoTable[216] = {4'b0000, 6'b100011, readAbsY, aluInT, aluCmp};
InfoTable[217] = {4'b0000, 6'b000000, push, aluInX, aluInp};
InfoTable[218] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[219] = {4'b0000, 6'b000000, readAbs, aluInXXX, aluXXX};
InfoTable[220] = {4'b0000, 6'b100011, readAbsX, aluInT, aluCmp};
InfoTable[221] = {4'b0000, 6'b100010, rmwAbsX, aluInT, aluDec};
InfoTable[222] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[223] = {4'b0000, 6'b100011, immediate, aluInT, aluCpx};
InfoTable[224] = {4'b1000, 6'b110011, readIndX, aluInT, aluSbc};
InfoTable[225] = {4'b0000, 6'b000000, immediate, aluInXXX, aluXXX};
InfoTable[226] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[227] = {4'b0000, 6'b100011, readZp, aluInT, aluCpx};
InfoTable[228] = {4'b1000, 6'b110011, readZp, aluInT, aluSbc};
InfoTable[229] = {4'b0000, 6'b100010, rmwZp, aluInT, aluInc};
InfoTable[230] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[231] = {4'b0100, 6'b100010, implied, aluInX, aluInc};
InfoTable[232] = {4'b1000, 6'b110011, immediate, aluInT, aluSbc};
InfoTable[233] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[234] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[235] = {4'b0000, 6'b100011, readAbs, aluInT, aluCpx};
InfoTable[236] = {4'b1000, 6'b110011, readAbs, aluInT, aluSbc};
InfoTable[237] = {4'b0000, 6'b100010, rmwAbs, aluInT, aluInc};
InfoTable[238] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[239] = {4'b0000, 6'b000000, relative, aluInXXX, aluXXX};
InfoTable[240] = {4'b1000, 6'b110011, readIndY, aluInT, aluSbc};
InfoTable[241] = {4'b1000, 6'b110011, readInd, aluInT, aluSbc};
InfoTable[242] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[243] = {4'b0000, 6'b000000, immediate, aluInXXX, aluXXX};
InfoTable[244] = {4'b1000, 6'b110011, readZpX, aluInT, aluSbc};
InfoTable[245] = {4'b0000, 6'b100010, rmwZpX, aluInT, aluInc};
InfoTable[246] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[247] = {4'b0000, 6'b001000, implied, aluInSet, aluXXX};
InfoTable[248] = {4'b1000, 6'b110011, readAbsY, aluInT, aluSbc};
InfoTable[249] = {4'b0100, 6'b100010, pop, aluInT, aluInp};
InfoTable[250] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
InfoTable[251] = {4'b0000, 6'b000000, readAbs, aluInXXX, aluXXX};
InfoTable[252] = {4'b1000, 6'b110011, readAbsX, aluInT, aluSbc};
InfoTable[253] = {4'b0000, 6'b100010, rmwAbsX, aluInT, aluInc};
InfoTable[254] = {4'b0000, 6'b000000, implied, aluInXXX, aluXXX};
end

    
    reg [0:43]       opcInfo;
    wire [0:43]      nextOpcInfo;		// Next  (decoded)
    wire [0:43]      nextOpcInfoReg;		// Next  (decoded) pipelined
    reg [7:0]        theOpcode;
    reg [7:0]        nextOpcode;
    
    // Program counter
    reg [15:0]       PC;		// Program counter
    
    // Address generation
    parameter [3:0]  nextAddrDef_nextAddrHold = 0,
                     nextAddrDef_nextAddrIncr = 1,
                     nextAddrDef_nextAddrIncrL = 2,
                     nextAddrDef_nextAddrIncrH = 3,
                     nextAddrDef_nextAddrDecrH = 4,
                     nextAddrDef_nextAddrPc = 5,
                     nextAddrDef_nextAddrIrq = 6,
                     nextAddrDef_nextAddrReset = 7,
                     nextAddrDef_nextAddrAbs = 8,
                     nextAddrDef_nextAddrAbsIndexed = 9,
                     nextAddrDef_nextAddrZeroPage = 10,
                     nextAddrDef_nextAddrZPIndexed = 11,
                     nextAddrDef_nextAddrStack = 12,
                     nextAddrDef_nextAddrRelative = 13;
    // Increment low bits only (zeropage accesses)
    // Increment high bits only (page-boundary)
    // Decrement high bits (branch backwards)
    reg [3:0]        nextAddr;
    reg [15:0]       myAddr;
    wire [15:0]      myAddrIncr;
    wire [7:0]       myAddrIncrH;
    wire [7:0]       myAddrDecrH;
    reg              theWe;
    reg              irqActive;
    // Output register
    reg [7:0]        doReg;
    // Buffer register
    reg [7:0]        T;
    // General registers
    reg [7:0]        A;		// Accumulator
    reg [7:0]        X;		// Index X
    reg [7:0]        Y;		// Index Y
    reg [7:0]        S;		// stack pointer
    // Status register
    reg              C;		// Carry
    reg              Z;		// Zero flag
    reg              I;		// Interrupt flag
    reg              D;		// Decimal mode
    wire             B;		// Break software interrupt
    reg              R;		// always 1
    reg              V;		// Overflow
    reg              N;		// Negative
    
    // ALU
    // ALU input
    reg [7:0]        aluInput;
    reg [7:0]        aluCmpInput;
    // ALU output
    reg [7:0]        aluRegisterOut;
    reg [7:0]        aluRmwOut;
    reg              aluC;
    reg              aluZ;
    reg              aluV;
    reg              aluN;
    // Indexing
    reg [8:0]        indexOut;
    
    wire             realbrk;
    
    always @(clk or opcInfo or A or X or Y or T or S)
    begin: processAluInput
        reg [7:0]        temp;
        temp = {8{1'b1}};
        
        if (opcInfo[opcInA] == 1'b1)
            temp = temp & A;
        if (opcInfo[opcInX] == 1'b1)
            temp = temp & X;
        if (opcInfo[opcInY] == 1'b1)
            temp = temp & Y;
        if (opcInfo[opcInS] == 1'b1)
            temp = temp & S;
        if (opcInfo[opcInT] == 1'b1)
            temp = temp & T;
        if (opcInfo[opcInBrk] == 1'b1)
            temp = temp & 8'b11100111;		// also DMB clear D (bit 3)
        if (opcInfo[opcInClear] == 1'b1)
            temp = {8{1'b0}};
        
        aluInput <= temp;
    end
    
    
    always @(clk or opcInfo or A or X or Y)
    begin: processCmpInput
        reg [7:0]        temp;
        temp = {8{1'b1}};
        if (opcInfo[opcInCmp] == 1'b1)
            temp = temp & A;
        if (opcInfo[opcInCpx] == 1'b1)
            temp = temp & X;
        if (opcInfo[opcInCpy] == 1'b1)
            temp = temp & Y;
        
        aluCmpInput <= temp;
    end
    
    // ALU consists of two parts
    // Read-Modify-Write or index instructions: INC/DEC/ASL/LSR/ROR/ROL 
    // Accumulator instructions: ADC, SBC, EOR, AND, EOR, ORA
    // Some instructions are both RMW and accumulator so for most
    // instructions the rmw results are routed through accu alu too.
    
    //	The B flag
    //----------
    //No actual "B" flag exists inside the 6502's processor status register. The B 
    //flag only exists in the status flag byte pushed to the stack. Naturally, 
    //when the flags are restored (via PLP or RTI), the B bit is discarded.
    //
    //Depending on the means, the B status flag will be pushed to the stack as 
    //either 0 or 1.
    //
    //software instructions BRK & PHP will push the B flag as being 1.
    //hardware interrupts IRQ & NMI will push the B flag as being 0.
    
function [7:0] trunc_to_8(input [31:0] val32);
  trunc_to_8 = val32[7:0];
endfunction

    always @(clk or opcInfo or aluInput or aluCmpInput or A or T or irqActive or N or V or R or D or I or Z or C)
    begin: processAlu
        reg [5:0]        lowBits;
        reg [8:0]        nineBits;
        reg [8:0]        rmwBits;
        reg [8:0]        tsxBits;
        
        reg              varC;
        reg              varZ;
        reg              varV;
        reg              varN;
        lowBits = {6{1'bx}};
        nineBits = {9{1'bx}};
        rmwBits = {9{1'bx}};
        tsxBits = {9{1'bx}};
        R <= 1'b1;
        
        // Shift unit
        case (opcInfo[aluMode1From:aluMode1To])
            aluModeInp :
                rmwBits = {C, aluInput};
            aluModeP :		// irqActive
                rmwBits = {C, N, V, R, ((~irqActive)), D, I, Z, C};
            aluModeInc :
                rmwBits = {C, trunc_to_8(aluInput +1)};
            aluModeDec :
                rmwBits = {C, trunc_to_8(aluInput - 1)};
            aluModeAsl :
                rmwBits = {aluInput, 1'b0};
            aluModeTSB :		// added by alan for 65c02
                begin
                    rmwBits = {1'b0, (aluInput[7:0] | A)};
                    tsxBits = {1'b0, (aluInput[7:0] & A)};
                end
            aluModeTRB :		// added by alan for 65c02
                begin
                    rmwBits = {1'b0, (aluInput[7:0] & ((~A)))};
                    tsxBits = {1'b0, (aluInput[7:0] & A)};
                end
            aluModeFlg :
                rmwBits = {aluInput[0], aluInput};
            aluModeLsr :
                rmwBits = {aluInput[0], 1'b0, aluInput[7:1]};
            aluModeRol :
                rmwBits = {aluInput, C};
            aluModeRor :
                rmwBits = {aluInput[0], C, aluInput[7:1]};
            default :
                rmwBits = {C, aluInput};
        endcase
        
        // ALU
        case (opcInfo[aluMode2From:aluMode2To])
            aluModeAdc :
                begin
                    lowBits = ({1'b0, A[3:0], rmwBits[8]}) + ({1'b0, rmwBits[3:0], 1'b1});
                    nineBits = ({1'b0, A}) + ({1'b0, rmwBits[7:0]}) + ({8'b00000000, rmwBits[8]});
                end
            aluModeSbc :
                begin
                    lowBits = ({1'b0, A[3:0], rmwBits[8]}) + ({1'b0, ((~rmwBits[3:0])), 1'b1});
                    nineBits = ({1'b0, A}) + ({1'b0, ((~rmwBits[7:0]))}) + ({8'b00000000, rmwBits[8]});
                end
            aluModeCmp :
                nineBits = ({1'b0, aluCmpInput}) + ({1'b0, ((~rmwBits[7:0]))}) + 9'b000000001;
            aluModeAnd :
                nineBits = {rmwBits[8], (A & rmwBits[7:0])};
            aluModeEor :
                nineBits = {rmwBits[8], (A ^ rmwBits[7:0])};
            aluModeOra :
                nineBits = {rmwBits[8], (A | rmwBits[7:0])};
            aluModeNoF :
                nineBits = 9'b000110000;
            default :
                nineBits = rmwBits;
        endcase
        
        varV = aluInput[6];		// Default for BIT / PLP / RTI
        
        if (opcInfo[aluMode1From:aluMode1To] == aluModeFlg)
            varZ = rmwBits[1];
        else if ((opcInfo[aluMode1From:aluMode1To] == aluModeTSB) | (opcInfo[aluMode1From:aluMode1To] == aluModeTRB))
        begin
            if (tsxBits[7:0] == 8'h00)
                varZ = 1'b1;
            else
                varZ = 1'b0;
        end
        else if (nineBits[7:0] == 8'h00)
            varZ = 1'b1;
        else
            varZ = 1'b0;
        
        if ((opcInfo[aluMode1From:aluMode1To] == aluModeBit) | (opcInfo[aluMode1From:aluMode1To] == aluModeFlg))
            varN = rmwBits[7];
        else
            varN = nineBits[7];
        
        varC = nineBits[8];
        
        case (opcInfo[aluMode2From:aluMode2To])
            //		n Set if most significant bit of result is set; else cleared.
            //		v Set if signed overflow; cleared if valid signed result.
            //		z Set if result is zero; else cleared.
            //		c Set if unsigned overflow; cleared if valid unsigned result
            
            aluModeAdc :
                // decimal mode low bits correction, is done after setting Z flag.
                if (D == 1'b1)
                begin
                    if (lowBits[5:1] > 9)
                    begin
                        nineBits[3:0] = nineBits[3:0] + 6;
                        if (lowBits[5] == 1'b0)
                            nineBits[8:4] = nineBits[8:4] + 1;
                    end
                end
            default :
                ;
        endcase
        
        case (opcInfo[aluMode2From:aluMode2To])
            aluModeAdc :
                begin
                    // decimal mode high bits correction, is done after setting Z and N flags
                    varV = (A[7] ^ nineBits[7]) & (rmwBits[7] ^ nineBits[7]);
                    if (D == 1'b1)
                    begin
                        if (nineBits[8:4] > 9)
                        begin
                            nineBits[8:4] = nineBits[8:4] + 6;
                            varC = 1'b1;
                        end
                    end
                end
            
            aluModeSbc :
                begin
                    varV = (A[7] ^ nineBits[7]) & (((~rmwBits[7])) ^ nineBits[7]);
                    if (D == 1'b1)
                    begin
                        // Check for borrow (lower 4 bits)
                        if (lowBits[5] == 1'b0)
                            nineBits[7:0] = nineBits[7:0] - 6;
                        // Check for borrow (upper 4 bits)
                        if (nineBits[8] == 1'b0)
                            nineBits[8:4] = nineBits[8:4] - 6;
                    end
                end
            default :
                ;
        endcase
        
        // fix n and z flag for 65c02 adc sbc instructions in decimal mode
        case (opcInfo[aluMode2From:aluMode2To])
            aluModeAdc :
                if (D == 1'b1)
                begin
                    if (nineBits[7:0] == 8'h00)
                        varZ = 1'b1;
                    else
                        varZ = 1'b0;
                    varN = nineBits[7];
                end
            aluModeSbc :
                if (D == 1'b1)
                begin
                    if (nineBits[7:0] == 8'h00)
                        varZ = 1'b1;
                    else
                        varZ = 1'b0;
                    varN = nineBits[7];
                end
            default :
                ;
        endcase
        
        // DMB Remove Pipelining        		
        //	if rising_edge(clk) then	
        aluRmwOut <= rmwBits[7:0];
        aluRegisterOut <= nineBits[7:0];
        aluC <= varC;
        aluZ <= varZ;
        aluV <= varV;
        aluN <= varN;
    end
    //		end if;
    
    
    always @(posedge clk)
    begin: calcInterrupt
        
        begin
            if (enable == 1'b1)
            begin
                if (theCpuCycle == cpuCycles_cycleStack4 | reset == 1'b0)
                    nmiReg <= 1'b1;
                if (nextCpuCycle != cpuCycles_cycleBranchTaken & nextCpuCycle != cpuCycles_Fetch)
                begin
                    irqReg <= irq_n;
                    nmiEdge <= nmi_n;
                    if ((nmiEdge == 1'b1) & (nmi_n == 1'b0))
                        nmiReg <= 1'b0;
                end
                // The 'or opcInfo(opcSetI)' prevents NMI immediately after BRK or IRQ.
                // Presumably this is done in the real 6502/6510 to prevent a double IRQ.
                processIrq <= (~((nmiReg & (irqReg | I)) | opcInfo[opcIRQ]));
            end
        end
    end
    
    //pipeirq: process(clk)
    //	begin
    //		if rising_edge(clk) then
    //			if enable = '1' then
    //				if (reset = '0') or (theCpuCycle = Fetch) then
    //                    -- The 'or opcInfo(opcSetI)' prevents NMI immediately after BRK or IRQ.
    //                    -- Presumably this is done in the real 6502/6510 to prevent a double IRQ.
    //                    processIrq <= not ((nmiReg and (irqReg or I)) or opcInfo(opcIRQ));
    //				end if;
    //			end if;
    //		end if;
    //	end process;
    
    
    always @(clk or di or reset or processIrq)
    begin: calcNextOpcode
        reg [7:0]        myNextOpcode;
        // Next  is read from input unless a reset or IRQ is pending.
        myNextOpcode = di;
        
        if (reset == 1'b0)
            myNextOpcode = 8'h4C;
        else if (processIrq == 1'b1)
            myNextOpcode = 8'h00;
        nextOpcode <= myNextOpcode;
    end
    
    assign nextOpcInfo = InfoTable[nextOpcode];
    
    // DMB Remove Pipelining        		
    //	process(clk)
    //	begin
    //		if rising_edge(clk) then
    assign nextOpcInfoReg = nextOpcInfo;
    //		end if;
    //	end process;
    
    // Read bits and flags from InfoTable and store in opcInfo.
    // This info is used to control the execution of the .
    
    always @(posedge clk)
    begin: calcOpcInfo
        
        begin
            if (enable == 1'b1)
            begin
                if ((reset == 1'b0) | (theCpuCycle == cpuCycles_Fetch))
                    opcInfo <= nextOpcInfo;
            end
        end
    end
    
    
    always @(posedge clk)
    begin: calcTheOpcode
        
        begin
            if (enable == 1'b1)
            begin
                if (theCpuCycle == cpuCycles_Fetch)
                begin
                    irqActive <= 1'b0;
                    if (processIrq == 1'b1)
                        irqActive <= 1'b1;
                    // Fetch 
                    theOpcode <= nextOpcode;
                end
            end
        end
    end
    
    // -----------------------------------------------------------------------
    // State machine
    // -----------------------------------------------------------------------
    
    always @(enable or theCpuCycle or opcInfo)
    begin
        updateRegisters <= 1'b0;
        if (enable == 1'b1)
        begin
            if (opcInfo[opcRti] == 1'b1)
            begin
                if (theCpuCycle == cpuCycles_cycleRead)
                    updateRegisters <= 1'b1;
            end
            else if (theCpuCycle == cpuCycles_Fetch)
                updateRegisters <= 1'b1;
        end
    end
    
    
    always @(posedge clk)
        
        begin
            if (enable == 1'b1)
                theCpuCycle <= nextCpuCycle;
            if (reset == 1'b0)
                theCpuCycle <= cpuCycles_cycle2;
        end
    
    // Determine the next cpu cycle. After the last cycle we always
    // go to Fetch to get the next opcode.
    
    always @(theCpuCycle or opcInfo or theOpcode or indexOut or T or N or V or C or Z)
    begin: calcNextCpuCycle
        nextCpuCycle <= cpuCycles_Fetch;
        
        case (theCpuCycle)
            cpuCycles_Fetch :
                nextCpuCycle <= cpuCycles_cycle2;
            cpuCycles_cycle2 :
                if (opcInfo[opcBranch] == 1'b1)
                begin
                    if ((N == theOpcode[5] & theOpcode[7:6] == 2'b00) | (V == theOpcode[5] & theOpcode[7:6] == 2'b01) | (C == theOpcode[5] & theOpcode[7:6] == 2'b10) | (Z == theOpcode[5] & theOpcode[7:6] == 2'b11) | (theOpcode[7:0] == 8'h80))		// Branch condition is true
                        nextCpuCycle <= cpuCycles_cycleBranchTaken;
                end
                else if (opcInfo[opcStackUp] == 1'b1)
                    nextCpuCycle <= cpuCycles_cycleStack1;
                else if (opcInfo[opcStackAddr] == 1'b1 & opcInfo[opcStackData] == 1'b1)
                    nextCpuCycle <= cpuCycles_cycleStack2;
                else if (opcInfo[opcStackAddr] == 1'b1)
                    nextCpuCycle <= cpuCycles_cycleStack1;
                else if (opcInfo[opcStackData] == 1'b1)
                    nextCpuCycle <= cpuCycles_cycleWrite;
                else if (opcInfo[opcAbsolute] == 1'b1)
                    nextCpuCycle <= cpuCycles_cycle3;
                else if (opcInfo[opcIndirect] == 1'b1)
                begin
                    if (opcInfo[indexX] == 1'b1)
                        nextCpuCycle <= cpuCycles_cyclePreIndirect;
                    else
                        nextCpuCycle <= cpuCycles_cycleIndirect;
                end
                else if (opcInfo[opcZeroPage] == 1'b1)
                begin
                    if (opcInfo[opcWrite] == 1'b1)
                    begin
                        if ((opcInfo[indexX] == 1'b1) | (opcInfo[indexY] == 1'b1))
                            nextCpuCycle <= cpuCycles_cyclePreWrite;
                        else
                            nextCpuCycle <= cpuCycles_cycleWrite;
                    end
                    else
                        if ((opcInfo[indexX] == 1'b1) | (opcInfo[indexY] == 1'b1))
                            nextCpuCycle <= cpuCycles_cyclePreRead;
                        else
                            nextCpuCycle <= cpuCycles_cycleRead2;
                end
                else if (opcInfo[opcJump] == 1'b1)
                    nextCpuCycle <= cpuCycles_cycleJump;
            cpuCycles_cycle3 :
                begin
                    nextCpuCycle <= cpuCycles_cycleRead;
                    if (opcInfo[opcWrite] == 1'b1)
                    begin
                        if ((opcInfo[indexX] == 1'b1) | (opcInfo[indexY] == 1'b1))
                            nextCpuCycle <= cpuCycles_cyclePreWrite;
                        else
                            nextCpuCycle <= cpuCycles_cycleWrite;
                    end
                    if ((opcInfo[opcIndirect] == 1'b1) & (opcInfo[indexX] == 1'b1))
                    begin
                        if (opcInfo[opcWrite] == 1'b1)
                            nextCpuCycle <= cpuCycles_cycleWrite;
                        else
                            nextCpuCycle <= cpuCycles_cycleRead2;
                    end
                end
            cpuCycles_cyclePreIndirect :
                nextCpuCycle <= cpuCycles_cycleIndirect;
            cpuCycles_cycleIndirect :
                nextCpuCycle <= cpuCycles_cycle3;
            cpuCycles_cycleBranchTaken :
                if (indexOut[8] != T[7])
                    nextCpuCycle <= cpuCycles_cycleBranchPage;
            cpuCycles_cyclePreRead :
                if (opcInfo[opcZeroPage] == 1'b1)
                    nextCpuCycle <= cpuCycles_cycleRead2;
            cpuCycles_cycleRead :
                if (opcInfo[opcJump] == 1'b1)
                    nextCpuCycle <= cpuCycles_cycleJump;
                else if (indexOut[8] == 1'b1)
                    nextCpuCycle <= cpuCycles_cycleRead2;
                else if (opcInfo[opcRmw] == 1'b1)
                begin
                    nextCpuCycle <= cpuCycles_cycleRmw;
                    if (opcInfo[indexX] == 1'b1 | opcInfo[indexY] == 1'b1)
                        nextCpuCycle <= cpuCycles_cycleRead2;
                end
            cpuCycles_cycleRead2 :
                if (opcInfo[opcRmw] == 1'b1)
                    nextCpuCycle <= cpuCycles_cycleRmw;
            cpuCycles_cycleRmw :
                nextCpuCycle <= cpuCycles_cycleWrite;
            cpuCycles_cyclePreWrite :
                nextCpuCycle <= cpuCycles_cycleWrite;
            cpuCycles_cycleStack1 :
                begin
                    nextCpuCycle <= cpuCycles_cycleRead;
                    if (opcInfo[opcStackAddr] == 1'b1)
                        nextCpuCycle <= cpuCycles_cycleStack2;
                end
            cpuCycles_cycleStack2 :
                begin
                    nextCpuCycle <= cpuCycles_cycleStack3;
                    if (opcInfo[opcRti] == 1'b1)
                        nextCpuCycle <= cpuCycles_cycleRead;
                    if (opcInfo[opcStackData] == 1'b0 & opcInfo[opcStackUp] == 1'b1)
                        nextCpuCycle <= cpuCycles_cycleJump;
                end
            cpuCycles_cycleStack3 :
                begin
                    nextCpuCycle <= cpuCycles_cycleRead;
                    if (opcInfo[opcStackData] == 1'b0 | opcInfo[opcStackUp] == 1'b1)
                        nextCpuCycle <= cpuCycles_cycleJump;
                    else if (opcInfo[opcStackAddr] == 1'b1)
                        nextCpuCycle <= cpuCycles_cycleStack4;
                end
            cpuCycles_cycleStack4 :
                nextCpuCycle <= cpuCycles_cycleRead;
            cpuCycles_cycleJump :
                if (opcInfo[opcIncrAfter] == 1'b1)
                    nextCpuCycle <= cpuCycles_cycleEnd;
            default :
                ;
        endcase
    end
    
    // -----------------------------------------------------------------------
    // T register
    // -----------------------------------------------------------------------
    
    always @(posedge clk)
    begin: calcT
        
        begin
            if (enable == 1'b1)
                case (theCpuCycle)
                    cpuCycles_cycle2 :
                        T <= di;
                    cpuCycles_cycleStack1, cpuCycles_cycleStack2 :
                        if (opcInfo[opcStackUp] == 1'b1)
                        begin
                            if (theOpcode == 8'h28 | theOpcode == 8'h40)		// plp or rti pulling the flags off the stack
                                T <= (di | 8'b00110000);		// Read from stack
                            else
                                T <= di;
                        end
                    cpuCycles_cycleIndirect, cpuCycles_cycleRead, cpuCycles_cycleRead2 :
                        T <= di;
                    default :
                        ;
                endcase
        end
    end
    
    // -----------------------------------------------------------------------
    // A register
    // -----------------------------------------------------------------------
    
    always @(posedge clk)
        
        begin
            if (updateRegisters)
            begin
                if (opcInfo[opcUpdateA] == 1'b1)
                    A <= aluRegisterOut;
            end
        end
    
    // -----------------------------------------------------------------------
    // X register
    // -----------------------------------------------------------------------
    
    always @(posedge clk)
        
        begin
            if (updateRegisters)
            begin
                if (opcInfo[opcUpdateX] == 1'b1)
                    X <= aluRegisterOut;
            end
        end
    
    // -----------------------------------------------------------------------
    // Y register
    // -----------------------------------------------------------------------
    
    always @(posedge clk)
        
        begin
            if (updateRegisters)
            begin
                if (opcInfo[opcUpdateY] == 1'b1)
                    Y <= aluRegisterOut;
            end
        end
    
    // -----------------------------------------------------------------------
    // C flag
    // -----------------------------------------------------------------------
    
    always @(posedge clk)
        
        begin
            if (updateRegisters)
            begin
                if (opcInfo[opcUpdateC] == 1'b1)
                    C <= aluC;
            end
        end
    
    // -----------------------------------------------------------------------
    // Z flag
    // -----------------------------------------------------------------------
    
    always @(posedge clk)
        
        begin
            if (updateRegisters)
            begin
                if (opcInfo[opcUpdateZ] == 1'b1)
                    Z <= aluZ;
            end
        end
    
    // -----------------------------------------------------------------------
    // I flag interupt flag
    // -----------------------------------------------------------------------
    
    always @(posedge clk or negedge reset)
        if (reset == 1'b0)
            I <= 1'b1;
        else 
        begin
            if (updateRegisters)
            begin
                if (opcInfo[opcUpdateI] == 1'b1)
                    I <= aluInput[2];
            end
        end
    // -----------------------------------------------------------------------
    // D flag
    // -----------------------------------------------------------------------
    
    always @(posedge clk or negedge reset)
        if (reset == 1'b0)
            D <= 1'b0;
        else 
        begin
            if (updateRegisters)
            begin
                if (opcInfo[opcUpdateD] == 1'b1)
                    D <= aluInput[3];
            end
        end
    
    // -----------------------------------------------------------------------
    // V flag
    // -----------------------------------------------------------------------
    
    always @(posedge clk)
        
        begin
            if (updateRegisters)
            begin
                if (opcInfo[opcUpdateV] == 1'b1)
                    V <= aluV;
            end
        end
    
    // -----------------------------------------------------------------------
    // N flag
    // -----------------------------------------------------------------------
    
    always @(posedge clk)
        
        begin
            if (updateRegisters)
            begin
                if (opcInfo[opcUpdateN] == 1'b1)
                    N <= aluN;
            end
        end
    
    // -----------------------------------------------------------------------
    // Stack pointer
    // -----------------------------------------------------------------------
    
    always @(posedge clk)
    begin: xhdl0
        reg [7:0]        sIncDec;
        reg              updateFlag;
        
        begin
            
            if (opcInfo[opcStackUp] == 1'b1)
                sIncDec = S + 1;
            else
                sIncDec = S - 1;
            
            if (enable == 1'b1)
            begin
                updateFlag = 1'b0;
                case (nextCpuCycle)
                    cpuCycles_cycleStack1 :
                        if ((opcInfo[opcStackUp] == 1'b1) | (opcInfo[opcStackData] == 1'b1))
                            updateFlag = 1'b1;
                    
                    cpuCycles_cycleStack2 :
                        updateFlag = 1'b1;
                    cpuCycles_cycleStack3 :
                        updateFlag = 1'b1;
                    cpuCycles_cycleStack4 :
                        updateFlag = 1'b1;
                    cpuCycles_cycleRead :
                        if (opcInfo[opcRti] == 1'b1)
                            updateFlag = 1'b1;
                    cpuCycles_cycleWrite :
                        if (opcInfo[opcStackData] == 1'b1)
                            updateFlag = 1'b1;
                    default :
                        ;
                endcase
                
                if (updateFlag)
                    S <= sIncDec;
            end
            
            if (updateRegisters)
            begin
                if (opcInfo[opcUpdateS] == 1'b1)
                    S <= aluRegisterOut;
            end
        end
    end
    
    // -----------------------------------------------------------------------
    // Data out
    // -----------------------------------------------------------------------
    
    always @(posedge clk)
    begin: calcDo
        
        begin
            if (enable == 1'b1)
            begin
                doReg <= aluRmwOut;
                case (nextCpuCycle)
                    cpuCycles_cycleStack2 :
                        if (opcInfo[opcIRQ] == 1'b1 & irqActive == 1'b0)
                            doReg <= myAddrIncr[15:8];
                        else
                            doReg <= PC[15:8];
                    cpuCycles_cycleStack3 :
                        doReg <= PC[7:0];
                    cpuCycles_cycleRmw :		// Read-modify-write write old value first.
                        doReg <= di;
                    default :
                        ;
                endcase
            end
        end
    end
    assign dout = doReg;
    
    // -----------------------------------------------------------------------
    // Write enable
    // -----------------------------------------------------------------------
    
    always @(posedge clk)
    begin: calcWe
        
        begin
            if (enable == 1'b1)
            begin
                theWe <= 1'b1;
                case (nextCpuCycle)
                    cpuCycles_cycleStack1 :
                        if (opcInfo[opcStackUp] == 1'b0 & ((opcInfo[opcStackAddr] == 1'b0) | (opcInfo[opcStackData] == 1'b1)))
                            theWe <= 1'b0;
                    cpuCycles_cycleStack2, cpuCycles_cycleStack3, cpuCycles_cycleStack4 :
                        if (opcInfo[opcStackUp] == 1'b0)
                            theWe <= 1'b0;
                    cpuCycles_cycleRmw :
                        theWe <= 1'b0;
                    cpuCycles_cycleWrite :
                        theWe <= 1'b0;
                    default :
                        ;
                endcase
            end
        end
    end
    //nwe <= theWe;
    assign nwe = theWe;
    
    // -----------------------------------------------------------------------
    // Program counter
    // -----------------------------------------------------------------------
    
    always @(posedge clk)
    begin: calcPC
        
        begin
            if (enable == 1'b1)
                case (theCpuCycle)
                    cpuCycles_Fetch :
                        PC <= myAddr;
                    cpuCycles_cycle2 :
                        if (irqActive == 1'b0)
                        begin
                            if (opcInfo[opcSecondByte] == 1'b1)
                                PC <= myAddrIncr;
                            else
                                PC <= myAddr;
                        end
                    cpuCycles_cycle3 :
                        if (opcInfo[opcAbsolute] == 1'b1)
                            PC <= myAddrIncr;
                    default :
                        ;
                endcase
        end
    end
    
    // -----------------------------------------------------------------------
    // Address generation
    // -----------------------------------------------------------------------
    
    always @(theCpuCycle or opcInfo or indexOut or T or reset)
    begin: calcNextAddr
        nextAddr <= nextAddrDef_nextAddrIncr;
        case (theCpuCycle)
            cpuCycles_cycle2 :
                if (opcInfo[opcStackAddr] == 1'b1 | opcInfo[opcStackData] == 1'b1)
                    nextAddr <= nextAddrDef_nextAddrStack;
                else if (opcInfo[opcAbsolute] == 1'b1)
                    nextAddr <= nextAddrDef_nextAddrIncr;
                else if (opcInfo[opcZeroPage] == 1'b1)
                    nextAddr <= nextAddrDef_nextAddrZeroPage;
                else if (opcInfo[opcIndirect] == 1'b1)
                    nextAddr <= nextAddrDef_nextAddrZeroPage;
                else if (opcInfo[opcSecondByte] == 1'b1)
                    nextAddr <= nextAddrDef_nextAddrIncr;
                else
                    nextAddr <= nextAddrDef_nextAddrHold;
            cpuCycles_cycle3 :
                if ((opcInfo[opcIndirect] == 1'b1) & (opcInfo[indexX] == 1'b1))
                    nextAddr <= nextAddrDef_nextAddrAbs;
                else
                    nextAddr <= nextAddrDef_nextAddrAbsIndexed;
            cpuCycles_cyclePreIndirect :
                nextAddr <= nextAddrDef_nextAddrZPIndexed;
            cpuCycles_cycleIndirect :
                nextAddr <= nextAddrDef_nextAddrIncrL;
            cpuCycles_cycleBranchTaken :
                nextAddr <= nextAddrDef_nextAddrRelative;
            cpuCycles_cycleBranchPage :
                if (T[7] == 1'b0)
                    nextAddr <= nextAddrDef_nextAddrIncrH;
                else
                    nextAddr <= nextAddrDef_nextAddrDecrH;
            cpuCycles_cyclePreRead :
                nextAddr <= nextAddrDef_nextAddrZPIndexed;
            cpuCycles_cycleRead :
                begin
                    nextAddr <= nextAddrDef_nextAddrPc;
                    if (opcInfo[opcJump] == 1'b1)
                        // Emulate 6510 bug, jmp(xxFF) fetches from same page.
                        // Replace with nextAddrIncr if emulating 65C02 or later cpu.
                        nextAddr <= nextAddrDef_nextAddrIncr;
                    //nextAddr <= nextAddrIncrL;	
                    else if (indexOut[8] == 1'b1)
                        nextAddr <= nextAddrDef_nextAddrIncrH;
                    else if (opcInfo[opcRmw] == 1'b1)
                        nextAddr <= nextAddrDef_nextAddrHold;
                end
            cpuCycles_cycleRead2 :
                begin
                    nextAddr <= nextAddrDef_nextAddrPc;
                    if (opcInfo[opcRmw] == 1'b1)
                        nextAddr <= nextAddrDef_nextAddrHold;
                end
            cpuCycles_cycleRmw :
                nextAddr <= nextAddrDef_nextAddrHold;
            cpuCycles_cyclePreWrite :
                begin
                    nextAddr <= nextAddrDef_nextAddrHold;
                    if (opcInfo[opcZeroPage] == 1'b1)
                        nextAddr <= nextAddrDef_nextAddrZPIndexed;
                    else if (indexOut[8] == 1'b1)
                        nextAddr <= nextAddrDef_nextAddrIncrH;
                end
            cpuCycles_cycleWrite :
                nextAddr <= nextAddrDef_nextAddrPc;
            cpuCycles_cycleStack1 :
                nextAddr <= nextAddrDef_nextAddrStack;
            cpuCycles_cycleStack2 :
                nextAddr <= nextAddrDef_nextAddrStack;
            cpuCycles_cycleStack3 :
                begin
                    nextAddr <= nextAddrDef_nextAddrStack;
                    if (opcInfo[opcStackData] == 1'b0)
                        nextAddr <= nextAddrDef_nextAddrPc;
                end
            cpuCycles_cycleStack4 :
                nextAddr <= nextAddrDef_nextAddrIrq;
            cpuCycles_cycleJump :
                nextAddr <= nextAddrDef_nextAddrAbs;
            
            default :
                ;
        endcase
        
        if (reset == 1'b0)
            nextAddr <= nextAddrDef_nextAddrReset;
    end
    
    
    always @(opcInfo or myAddr or T or X or Y)
    begin: indexAlu
        if (opcInfo[indexX] == 1'b1)
            indexOut <= ({1'b0, T}) + ({1'b0, X});
        else if (opcInfo[indexY] == 1'b1)
            indexOut <= ({1'b0, T}) + ({1'b0, Y});
        else if (opcInfo[opcBranch] == 1'b1)
            indexOut <= ({1'b0, T}) + ({1'b0, myAddr[7:0]});
        else
            indexOut <= {1'b0, T};
    end
    
    
    always @(posedge clk)
    begin: calcAddr
        
        begin
            if (enable == 1'b1)
                case (nextAddr)
                    nextAddrDef_nextAddrIncr :
                        myAddr <= myAddrIncr;
                    nextAddrDef_nextAddrIncrL :
                        myAddr[7:0] <= myAddrIncr[7:0];
                    nextAddrDef_nextAddrIncrH :
                        myAddr[15:8] <= myAddrIncrH;
                    nextAddrDef_nextAddrDecrH :
                        myAddr[15:8] <= myAddrDecrH;
                    nextAddrDef_nextAddrPc :
                        myAddr <= PC;
                    nextAddrDef_nextAddrIrq :
                        begin
                            myAddr <= 16'hFFFE;
                            if (nmiReg == 1'b0)
                                myAddr <= 16'hFFFA;
                        end
                    nextAddrDef_nextAddrReset :
                        myAddr <= 16'hFFFC;
                    nextAddrDef_nextAddrAbs :
                        myAddr <= {di, T};
                    nextAddrDef_nextAddrAbsIndexed :		//myAddr <= di & indexOut(7 downto 0);
                        if (theOpcode == 8'h7C)
                            myAddr <= ({di, T}) + ({8'h00, X});
                        else
                            myAddr <= {di, indexOut[7:0]};
                    nextAddrDef_nextAddrZeroPage :
                        myAddr <= {8'b00000000, di};
                    nextAddrDef_nextAddrZPIndexed :
                        myAddr <= {8'b00000000, indexOut[7:0]};
                    nextAddrDef_nextAddrStack :
                        myAddr <= {8'b00000001, S};
                    nextAddrDef_nextAddrRelative :
                        myAddr[7:0] <= indexOut[7:0];
                    default :
                        ;
                endcase
        end
    end
    
    assign myAddrIncr = myAddr + 1;
    assign myAddrIncrH = myAddr[15:8] + 1;
    assign myAddrDecrH = myAddr[15:8] - 1;
    assign addr = myAddr;
    
    // DMB This looked plain broken and inferred a latch
    //    
    //	calcsync: process(clk)
    //	begin
    //		
    //			if enable = '1' then
    //				case theCpuCycle is
    //				when Fetch =>			sync <= '1';
    //				when others =>					sync <= '0';			
    //				end case;
    //			end if;
    //	end process;
    
    assign sync = (theCpuCycle == cpuCycles_Fetch) ? 1'b1 : 
                  1'b0;
    
    assign sync_irq = irqActive;
    
    assign Regs = {PC, 8'b00000001, S, N, V, R, B, D, I, Z, C, Y, X, A};
    
endmodule


