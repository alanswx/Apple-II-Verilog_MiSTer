module R65C02
  (input  reset,
   input  clk,
   input  enable,
   input  nmi_n,
   input  irq_n,
   input  [7:0] di,
   output [7:0] dout,
   output [15:0] addr,
   output nwe,
   output sync,
   output sync_irq,
   output [63:0] Regs);
  wire [4:0] thecpucycle;
  wire [4:0] nextcpucycle;
  wire updateregisters;
  wire processirq;
  wire nmireg;
  wire nmiedge;
  wire irqreg;
  wire [43:0] opcinfo;
  wire [43:0] nextopcinfo;
  wire [7:0] theopcode;
  wire [7:0] nextopcode;
  wire [15:0] pc;
  wire [3:0] nextaddr;
  wire [15:0] myaddr;
  wire [15:0] myaddrincr;
  wire [7:0] myaddrincrh;
  wire [7:0] myaddrdecrh;
  wire thewe;
  wire irqactive;
  wire [7:0] doreg;
  wire [7:0] t;
  wire [7:0] a;
  wire [7:0] x;
  wire [7:0] y;
  wire [7:0] s;
  wire c;
  wire z;
  wire i;
  wire d;
  wire b;
  wire r;
  wire v;
  wire n;
  wire [7:0] aluinput;
  wire [7:0] alucmpinput;
  wire [7:0] aluregisterout;
  wire [7:0] alurmwout;
  wire aluc;
  wire aluz;
  wire aluv;
  wire alun;
  wire [8:0] indexout;
  wire n8_o;
  wire [7:0] n10_o;
  wire [7:0] n12_o;
  wire n14_o;
  wire [7:0] n15_o;
  wire [7:0] n16_o;
  wire n17_o;
  wire [7:0] n18_o;
  wire [7:0] n19_o;
  wire n20_o;
  wire [7:0] n21_o;
  wire [7:0] n22_o;
  wire n23_o;
  wire [7:0] n24_o;
  wire [7:0] n25_o;
  wire n26_o;
  wire [7:0] n28_o;
  wire [7:0] n29_o;
  wire n30_o;
  wire [7:0] n32_o;
  wire n37_o;
  wire [7:0] n39_o;
  wire [7:0] n41_o;
  wire n43_o;
  wire [7:0] n44_o;
  wire [7:0] n45_o;
  wire n46_o;
  wire [7:0] n47_o;
  wire [7:0] n48_o;
  wire [3:0] n60_o;
  wire [8:0] n61_o;
  wire n63_o;
  wire [1:0] n64_o;
  wire [2:0] n65_o;
  wire [3:0] n66_o;
  wire n67_o;
  wire [4:0] n68_o;
  wire [5:0] n69_o;
  wire [6:0] n70_o;
  wire [7:0] n71_o;
  wire [8:0] n72_o;
  wire n74_o;
  wire [7:0] n76_o;
  wire [8:0] n77_o;
  wire n79_o;
  wire [7:0] n81_o;
  wire [8:0] n82_o;
  wire n84_o;
  wire [8:0] n86_o;
  wire n88_o;
  wire [7:0] n89_o;
  wire [8:0] n91_o;
  wire [7:0] n92_o;
  wire [8:0] n94_o;
  wire n96_o;
  wire [7:0] n97_o;
  wire [7:0] n98_o;
  wire [8:0] n100_o;
  wire [7:0] n101_o;
  wire [8:0] n103_o;
  wire n105_o;
  wire n106_o;
  wire [8:0] n107_o;
  wire n109_o;
  wire n110_o;
  wire [1:0] n112_o;
  wire [6:0] n113_o;
  wire [8:0] n114_o;
  wire n116_o;
  wire [8:0] n117_o;
  wire n119_o;
  wire n120_o;
  wire [1:0] n121_o;
  wire [6:0] n122_o;
  wire [8:0] n123_o;
  wire n125_o;
  wire [8:0] n126_o;
  wire [10:0] n127_o;
  reg [8:0] n128_o;
  reg [8:0] n131_o;
  wire [2:0] n133_o;
  wire [3:0] n134_o;
  wire [4:0] n136_o;
  wire n137_o;
  wire [5:0] n138_o;
  wire [3:0] n139_o;
  wire [4:0] n141_o;
  wire [5:0] n143_o;
  wire [5:0] n144_o;
  wire [8:0] n146_o;
  wire [7:0] n147_o;
  wire [8:0] n149_o;
  wire [8:0] n150_o;
  wire n151_o;
  wire [8:0] n153_o;
  wire [8:0] n154_o;
  wire n156_o;
  wire [3:0] n157_o;
  wire [4:0] n159_o;
  wire n160_o;
  wire [5:0] n161_o;
  wire [3:0] n162_o;
  wire [3:0] n163_o;
  wire [4:0] n165_o;
  wire [5:0] n167_o;
  wire [5:0] n168_o;
  wire [8:0] n170_o;
  wire [7:0] n171_o;
  wire [7:0] n172_o;
  wire [8:0] n174_o;
  wire [8:0] n175_o;
  wire n176_o;
  wire [8:0] n178_o;
  wire [8:0] n179_o;
  wire n181_o;
  wire [8:0] n183_o;
  wire [7:0] n184_o;
  wire [7:0] n185_o;
  wire [8:0] n187_o;
  wire [8:0] n188_o;
  wire [8:0] n190_o;
  wire n192_o;
  wire n193_o;
  wire [7:0] n194_o;
  wire [7:0] n195_o;
  wire [8:0] n196_o;
  wire n198_o;
  wire n199_o;
  wire [7:0] n200_o;
  wire [7:0] n201_o;
  wire [8:0] n202_o;
  wire n204_o;
  wire n205_o;
  wire [7:0] n206_o;
  wire [7:0] n207_o;
  wire [8:0] n208_o;
  wire n210_o;
  wire n212_o;
  wire [6:0] n213_o;
  reg [5:0] n215_o;
  reg [8:0] n218_o;
  wire n220_o;
  wire [3:0] n221_o;
  wire n223_o;
  wire n224_o;
  wire [3:0] n225_o;
  wire n227_o;
  wire [3:0] n228_o;
  wire n230_o;
  wire n231_o;
  wire [7:0] n232_o;
  wire n234_o;
  wire n237_o;
  wire [7:0] n238_o;
  wire n240_o;
  wire n243_o;
  wire n244_o;
  wire n245_o;
  wire [3:0] n246_o;
  wire n248_o;
  wire [3:0] n249_o;
  wire n251_o;
  wire n252_o;
  wire n253_o;
  wire n254_o;
  wire n255_o;
  wire n256_o;
  wire [2:0] n257_o;
  wire [4:0] n258_o;
  wire n260_o;
  wire [3:0] n261_o;
  wire [3:0] n263_o;
  wire n264_o;
  wire n265_o;
  wire [4:0] n266_o;
  wire [8:0] n267_o;
  wire [4:0] n268_o;
  wire [4:0] n270_o;
  wire [4:0] n271_o;
  wire [4:0] n272_o;
  wire [8:0] n273_o;
  wire [8:0] n274_o;
  wire n275_o;
  wire n277_o;
  reg [8:0] n278_o;
  wire [2:0] n279_o;
  wire n280_o;
  wire n281_o;
  wire n282_o;
  wire n283_o;
  wire n284_o;
  wire n285_o;
  wire n286_o;
  wire [4:0] n287_o;
  wire n289_o;
  wire [4:0] n290_o;
  wire [4:0] n292_o;
  wire [4:0] n293_o;
  wire [4:0] n294_o;
  wire n296_o;
  wire n298_o;
  wire n299_o;
  wire n301_o;
  wire n302_o;
  wire n303_o;
  wire n304_o;
  wire n305_o;
  wire n306_o;
  wire n307_o;
  wire n308_o;
  wire n309_o;
  wire n310_o;
  wire n311_o;
  wire [7:0] n312_o;
  wire [7:0] n314_o;
  wire [7:0] n315_o;
  wire [7:0] n316_o;
  wire n317_o;
  wire [8:0] n318_o;
  wire n319_o;
  wire n320_o;
  wire n321_o;
  wire [8:0] n322_o;
  wire [4:0] n323_o;
  wire [4:0] n325_o;
  wire [3:0] n326_o;
  wire [3:0] n327_o;
  wire [3:0] n328_o;
  wire n329_o;
  wire [4:0] n330_o;
  wire [4:0] n331_o;
  wire [3:0] n332_o;
  wire [3:0] n333_o;
  wire [3:0] n334_o;
  wire [8:0] n335_o;
  wire [8:0] n336_o;
  wire n338_o;
  wire [1:0] n339_o;
  wire [3:0] n340_o;
  wire [3:0] n341_o;
  reg [3:0] n342_o;
  wire [4:0] n343_o;
  wire [4:0] n344_o;
  reg [4:0] n345_o;
  reg n347_o;
  reg n348_o;
  wire [2:0] n349_o;
  wire [8:0] n350_o;
  wire [7:0] n351_o;
  wire n353_o;
  wire n356_o;
  wire [8:0] n357_o;
  wire n358_o;
  wire n359_o;
  wire n360_o;
  wire n362_o;
  wire [8:0] n363_o;
  wire [7:0] n364_o;
  wire n366_o;
  wire n369_o;
  wire [8:0] n370_o;
  wire n371_o;
  wire n372_o;
  wire n373_o;
  wire n375_o;
  wire [1:0] n376_o;
  reg n377_o;
  reg n378_o;
  wire [7:0] n379_o;
  wire [8:0] n380_o;
  wire [7:0] n381_o;
  wire n388_o;
  wire n389_o;
  wire n390_o;
  wire n392_o;
  wire n394_o;
  wire n396_o;
  wire n397_o;
  wire n398_o;
  wire n399_o;
  wire n401_o;
  wire n402_o;
  wire n405_o;
  wire n406_o;
  wire n407_o;
  wire n408_o;
  wire n409_o;
  wire n412_o;
  wire n413_o;
  wire n419_o;
  reg n420_q;
  wire n421_o;
  reg n422_q;
  wire n423_o;
  reg n424_q;
  wire n425_o;
  reg n426_q;
  wire n429_o;
  wire [7:0] n431_o;
  wire [7:0] n433_o;
  wire [7:0] n438_o;
  localparam [11263:0] n440_o = "00000011001000111000000001010000000001000XXX10001000101001000010000000000001000000101XXX00000000001000000000000000XXXXXXXXXXXXXXXXXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000101010000000001000000001001100000XXX10001000101010000000000000000001000000101XXX00001000111010000000001000000001001010000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000000000010000000000XXXXXXXX0001000XXX10001000101000000000000000000001000000101XXX10001000110000000000000000100000001010000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000101100000000001000000001001100000XXX10001000101100000000000000000001000000101XXX00001000111100000000001000000001001010000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000001000000100000000XXXXXXXXXXXXXXXXXX10001000101001000001000000000001000000101XXX10001000101001000000000000000001000000101XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000101010000000001000000001001101000XXX10001000101010000010000000000001000000101XXX00001000111010000010001000000001001010000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000010000000000000000000000010100000XXX10001000101100000001000000000001000000101XXX10001000100000000000000000100000000010000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000101100000000001000000001001101000XXX10001000101100000010000000000001000000101XXX00001000111100000010001000000001001010000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000001000101000000000XXXXXXXXXXXXXXXXXX10001000101001000010000000000001000000100XXX00000000001000000000000000XXXXXXXXXXXXXXXXXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00001100101010000000000000000001000101100XXX10001000101010000000000000000001000000100XXX00001000111010000000001000000001001011000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00001111110000010000100000000001000100000XXX10001000101000000000000000000001000000100XXX10001000110000000000000000100000001011000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00001100101100000000000000000001000101100XXX10001000101100000000000000000001000000100XXX00001000111100000000001000000001001011000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000001000000100000000XXXXXXXXXXXXXXXXXX10001000101001000001000000000001000000100XXX10001000101001000000000000000001000000100XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00001100101010000010000000000001000101100XXX10001000101010000010000000000001000000100XXX00001000111010000010001000000001001011000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000010000000000000000000000000100000XXX10001000101100000001000000000001000000100XXX10001000100000000000000000100000000011000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00001100101100000010000000000001000101100XXX10001000101100000010000000000001000000100XXX00001000111100000010001000000001001011000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00001111110000111000100010000001000100000XXX10001000101001000010000000000001000000110XXX00000000001000000000000000XXXXXXXXXXXXXXXXXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000001000000000000000XXXXXXXXXXXXXXXXXX10001000101010000000000000000001000000110XXX00001000111010000000001000000001001000000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000000000010000000000100000000000000XXX10001000101000000000000000000001000000110XXX10001000110000000000000000100000001000000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000001000001000000000XXXXXXXXXXXXXXXXXX10001000101100000000000000000001000000110XXX00001000111100000000001000000001001000000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000001000000100000000XXXXXXXXXXXXXXXXXX10001000101001000001000000000001000000110XXX10001000101001000000000000000001000000110XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000001000000000000000XXXXXXXXXXXXXXXXXX10001000101010000010000000000001000000110XXX00001000111010000010001000000001001000000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX0000000100000000000000000000000001XXXXXXXXXX10001000101100000001000000000001000000110XXX00000000000000010000000000000100000000000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000001100000000000000XXXXXXXXXXXXXXXXXX10001000101100000010000000000001000000110XXX00001000111100000010001000000001001000000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000000000101000100100XXXXXXXXXXXXXXXXXX10001100111001000010000000000001000000010XXX00000000001000000000000000XXXXXXXXXXXXXXXXXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000001010000000010000000000010000000XXX10001100111010000000000000000001000000010XXX00001000111010000000001000000001001001000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX10001000100000010000100000000001000000000XXX10001100111000000000000000000001000000010XXX10001000110000000000000000100000001001000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000001100001000000000XXXXXXXXXXXXXXXXXX10001100111100000000000000000001000000010XXX00001000111100000000001000000001001001000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000001000000100000000XXXXXXXXXXXXXXXXXX10001100111001000001000000000001000000010XXX10001100111001000000000000000001000000010XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000001010000010010000000000010000000XXX10001100111010000010000000000001000000010XXX00001000111010000010001000000001001001000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX0000000100000000000000000000000000XXXXXXXXXX10001100111100000001000000000001000000010XXX00101000100000010000100000000001000000000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000001100001010000000XXXXXXXXXXXXXXXXXX10001100111100000010000000000001000000010XXX00001000111100000010001000000001001001000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000001000000100000000XXXXXXXXXXXXXXXXXX00000000001001000010010000100000000000000XXX00000000001000000000000000XXXXXXXXXXXXXXXXXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000001010000000010000000100000000000XXX00000000001010000000010000100000000000000XXX00000000001010000000010000001000000000000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00101000100000000000000000000100000011000XXX00000000101000000000000000000001000101100XXX10001000100000000000000000001000000000000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000001100000000010000000100000000000XXX00000000001100000000010000100000000000000XXX00000000001100000000010000001000000000000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000001000000100000000XXXXXXXXXXXXXXXXXX00000000001001000001010000100000000000000XXX00000000001001000000010000100000000000000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000001010000010010000000100000000000XXX00000000001010000010010000100000000000000XXX00000000001010000001010000001000000000000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX10001000100000000000000000000100000000000XXX00000000001100000001010000100000000000000XXX00010000000000000000000000001000000000000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000001100000000010000000000010000000XXX00000000001100000010010000100000000000000XXX00000000001100000010010000000000010000000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00101000101000000000000000000001000000000XXX10001000101001000010000000000001000000000XXX01001000101000000000000000000001000000000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00101000101010000000000000000001000000000XXX10001000101010000000000000000001000000000XXX01001000101010000000000000000001000000000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00101000100000000000000000100000000000000XXX10001000101000000000000000000001000000000XXX01001000100000000000000000100000000000000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00101000101100000000000000000001000000000XXX10001000101100000000000000000001000000000XXX01001000101100000000000000000001000000000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000001000000100000000XXXXXXXXXXXXXXXXXX10001000101001000001000000000001000000000XXX10001000101001000000000000000001000000000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00101000101010000010000000000001000000000XXX10001000101010000010000000000001000000000XXX01001000101010000001000000000001000000000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000100000000000000000000000000010100000XXX10001000101100000001000000000001000000000XXX01001000100000000000000000000010000000000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00101000101100000010000000000001000000000XXX10001000101100000010000000000001000000000XXX01001000101100000001000000000001000000000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX000010001110000000000000000000010000000010010000100011100100001000000000000100000000110000000000001000000000000000XXXXXXXXXXXXXXXXXX00000000000000000000000000XXXXXXXXXXXXXXXXXX000010001110100000000000000000010000000010010000100011101000000000000000000100000000110000001000101010000000001000000001000011000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00101000100000000000000000000100000010000XXX0000100011100000000000000000000100000000110001001000100000000000000000001000000011000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX000010001111000000000000000000010000000010010000100011110000000000000000000100000000110000001000101100000000001000000001000011000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000001000000100000000XXXXXXXXXXXXXXXXXX000010001110010000010000000000010000000011000000100011100100000000000000000100000000110000000000000000000000000000XXXXXXXXXXXXXXXXXX00000000001000000000000000XXXXXXXXXXXXXXXXXX0000100011101000001000000000000100000000110000001000101010000010001000000001000011000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX0000001000000000000000000000000001XXXXXXXXXX0000100011110000000100000000000100000000110000000000000000010000000000001000000000000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000001100000000000000XXXXXXXXXXXXXXXXXX0000100011110000001000000000000100000000110000001000101100000010001000000001000011000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX0000100011100000000000000000000100000000101010001100111001000010000000000001000000011XXX00000000001000000000000000XXXXXXXXXXXXXXXXXX00000000000000000000000000XXXXXXXXXXXXXXXXXX0000100011101000000000000000000100000000101010001100111010000000000000000001000000011XXX00001000101010000000001000000001000010000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX01001000100000000000000000001000000010000XXX10001100111000000000000000000001000000011XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000000000000000000000XXXXXXXXXXXXXXXXXX0000100011110000000000000000000100000000101010001100111100000000000000000001000000011XXX00001000101100000000001000000001000010000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000001000000100000000XXXXXXXXXXXXXXXXXX10001100111001000001000000000001000000011XXX10001100111001000000000000000001000000011XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000001000000000000000XXXXXXXXXXXXXXXXXX10001100111010000010000000000001000000011XXX00001000101010000010001000000001000010000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX0000001000000000000000000000000000XXXXXXXXXX10001100111100000001000000000001000000011XXX01001000100000010000100000000001000000000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX00000000001100000000000000XXXXXXXXXXXXXXXXXX10001100111100000010000000000001000000011XXX00001000101100000010001000000001000010000XXX00000000000000000000000000XXXXXXXXXXXXXXXXXX";
  wire n444_o;
  wire n446_o;
  wire n447_o;
  wire n449_o;
  wire [43:0] n452_o;
  reg [43:0] n453_q;
  wire n457_o;
  wire n460_o;
  wire n464_o;
  wire n465_o;
  wire [7:0] n469_o;
  reg [7:0] n470_q;
  wire n471_o;
  reg n472_q;
  wire n475_o;
  wire n477_o;
  wire n480_o;
  wire n482_o;
  wire n485_o;
  wire n486_o;
  wire n488_o;
  wire [4:0] n494_o;
  wire n495_o;
  wire [4:0] n497_o;
  reg [4:0] n500_q;
  wire n503_o;
  wire n504_o;
  wire n505_o;
  wire n506_o;
  wire [1:0] n507_o;
  wire n509_o;
  wire n510_o;
  wire n511_o;
  wire n512_o;
  wire [1:0] n513_o;
  wire n515_o;
  wire n516_o;
  wire n517_o;
  wire n518_o;
  wire n519_o;
  wire [1:0] n520_o;
  wire n522_o;
  wire n523_o;
  wire n524_o;
  wire n525_o;
  wire n526_o;
  wire [1:0] n527_o;
  wire n529_o;
  wire n530_o;
  wire n531_o;
  wire n533_o;
  wire n534_o;
  wire [4:0] n537_o;
  wire n538_o;
  wire n539_o;
  wire n540_o;
  wire n541_o;
  wire n542_o;
  wire n543_o;
  wire n544_o;
  wire n545_o;
  wire n546_o;
  wire [4:0] n549_o;
  wire n550_o;
  wire n551_o;
  wire n552_o;
  wire n553_o;
  wire n554_o;
  wire [4:0] n557_o;
  wire n558_o;
  wire n559_o;
  wire n560_o;
  wire [4:0] n563_o;
  wire [4:0] n564_o;
  wire n565_o;
  wire [4:0] n568_o;
  wire [4:0] n569_o;
  wire [4:0] n570_o;
  wire [4:0] n572_o;
  wire [4:0] n574_o;
  wire [4:0] n576_o;
  wire [4:0] n578_o;
  wire [4:0] n580_o;
  wire [4:0] n581_o;
  wire n583_o;
  wire n584_o;
  wire n585_o;
  wire n586_o;
  wire n587_o;
  wire [4:0] n590_o;
  wire [4:0] n592_o;
  wire n594_o;
  wire n595_o;
  wire n596_o;
  wire n597_o;
  wire [4:0] n600_o;
  wire [4:0] n601_o;
  wire n603_o;
  wire n605_o;
  wire n607_o;
  wire n608_o;
  wire n609_o;
  wire n610_o;
  wire [4:0] n613_o;
  wire n615_o;
  wire n616_o;
  wire [4:0] n619_o;
  wire n621_o;
  wire n622_o;
  wire n623_o;
  wire n624_o;
  wire n625_o;
  wire n626_o;
  wire n627_o;
  wire [4:0] n630_o;
  wire [4:0] n633_o;
  wire [4:0] n635_o;
  wire [4:0] n637_o;
  wire n639_o;
  wire n640_o;
  wire [4:0] n643_o;
  wire n645_o;
  wire n647_o;
  wire n649_o;
  wire n650_o;
  wire [4:0] n653_o;
  wire n656_o;
  wire n657_o;
  wire [4:0] n660_o;
  wire n662_o;
  wire n663_o;
  wire n664_o;
  wire n665_o;
  wire [4:0] n667_o;
  wire n669_o;
  wire n670_o;
  wire n671_o;
  wire n672_o;
  wire n673_o;
  wire n674_o;
  wire [4:0] n677_o;
  wire [4:0] n679_o;
  wire n682_o;
  wire n684_o;
  wire n685_o;
  wire [4:0] n688_o;
  wire n690_o;
  wire [15:0] n691_o;
  reg [4:0] n699_o;
  wire n705_o;
  wire n706_o;
  wire n708_o;
  wire n710_o;
  wire n711_o;
  wire [7:0] n713_o;
  wire [7:0] n714_o;
  wire [7:0] n715_o;
  wire n717_o;
  wire n719_o;
  wire n720_o;
  wire n722_o;
  wire n724_o;
  wire n725_o;
  wire n727_o;
  wire n728_o;
  wire [2:0] n729_o;
  reg [7:0] n730_o;
  wire [7:0] n734_o;
  reg [7:0] n735_q;
  wire n739_o;
  wire n741_o;
  wire [7:0] n744_o;
  reg [7:0] n745_q;
  wire n749_o;
  wire n751_o;
  wire [7:0] n754_o;
  reg [7:0] n755_q;
  wire n759_o;
  wire n761_o;
  wire [7:0] n764_o;
  reg [7:0] n765_q;
  wire n769_o;
  wire n771_o;
  wire n774_o;
  reg n775_q;
  wire n779_o;
  wire n781_o;
  wire n784_o;
  reg n785_q;
  wire n788_o;
  wire n790_o;
  wire n791_o;
  wire n793_o;
  wire n798_o;
  reg n799_q;
  wire n802_o;
  wire n804_o;
  wire n805_o;
  wire n807_o;
  wire n812_o;
  reg n813_q;
  wire n817_o;
  wire n819_o;
  wire n822_o;
  reg n823_q;
  wire n827_o;
  wire n829_o;
  wire n832_o;
  reg n833_q;
  wire n839_o;
  wire [7:0] n841_o;
  wire [7:0] n843_o;
  wire [7:0] n844_o;
  wire n845_o;
  wire n846_o;
  wire n847_o;
  wire n850_o;
  wire n852_o;
  wire n854_o;
  wire n856_o;
  wire n858_o;
  wire n859_o;
  wire n862_o;
  wire n864_o;
  wire n865_o;
  wire n868_o;
  wire n870_o;
  wire [5:0] n871_o;
  reg n876_o;
  wire [7:0] n878_o;
  wire n879_o;
  wire n881_o;
  wire [7:0] n882_o;
  wire n883_o;
  reg [7:0] n888_q;
  wire n891_o;
  wire n892_o;
  wire n893_o;
  wire [7:0] n894_o;
  wire [7:0] n895_o;
  wire [7:0] n896_o;
  wire n898_o;
  wire [7:0] n899_o;
  wire n901_o;
  wire n903_o;
  wire [2:0] n904_o;
  reg [7:0] n905_o;
  wire [7:0] n909_o;
  reg [7:0] n910_q;
  wire n913_o;
  wire n914_o;
  wire n915_o;
  wire n916_o;
  wire n917_o;
  wire n918_o;
  wire n919_o;
  wire n922_o;
  wire n924_o;
  wire n925_o;
  wire n926_o;
  wire n929_o;
  wire n931_o;
  wire n933_o;
  wire n934_o;
  wire n936_o;
  wire n937_o;
  wire n939_o;
  wire n941_o;
  wire [3:0] n942_o;
  reg n946_o;
  wire n951_o;
  reg n952_q;
  wire n956_o;
  wire n957_o;
  wire n958_o;
  wire [15:0] n959_o;
  wire [15:0] n960_o;
  wire n962_o;
  wire n963_o;
  wire [15:0] n964_o;
  wire n966_o;
  wire [2:0] n967_o;
  reg [15:0] n968_o;
  wire [15:0] n972_o;
  reg [15:0] n973_q;
  wire n975_o;
  wire n976_o;
  wire n977_o;
  wire n978_o;
  wire n979_o;
  wire n980_o;
  wire n981_o;
  wire [3:0] n984_o;
  wire [3:0] n986_o;
  wire [3:0] n988_o;
  wire [3:0] n990_o;
  wire [3:0] n992_o;
  wire n994_o;
  wire n995_o;
  wire n996_o;
  wire n997_o;
  wire [3:0] n1000_o;
  wire n1002_o;
  wire n1004_o;
  wire n1006_o;
  wire n1008_o;
  wire n1009_o;
  wire n1010_o;
  wire [3:0] n1013_o;
  wire n1015_o;
  wire n1017_o;
  wire n1018_o;
  wire n1019_o;
  wire n1020_o;
  wire [3:0] n1023_o;
  wire [3:0] n1025_o;
  wire [3:0] n1027_o;
  wire n1030_o;
  wire n1031_o;
  wire [3:0] n1034_o;
  wire n1037_o;
  wire n1039_o;
  wire n1040_o;
  wire n1041_o;
  wire [3:0] n1044_o;
  wire [3:0] n1046_o;
  wire n1049_o;
  wire n1051_o;
  wire n1053_o;
  wire n1055_o;
  wire n1056_o;
  wire n1057_o;
  wire [3:0] n1060_o;
  wire n1063_o;
  wire n1065_o;
  wire n1067_o;
  wire [16:0] n1068_o;
  reg [3:0] n1080_o;
  wire n1082_o;
  wire [3:0] n1084_o;
  wire n1087_o;
  wire [8:0] n1089_o;
  wire [8:0] n1091_o;
  wire [8:0] n1092_o;
  wire n1093_o;
  wire [8:0] n1095_o;
  wire [8:0] n1097_o;
  wire [8:0] n1098_o;
  wire n1099_o;
  wire [8:0] n1101_o;
  wire [7:0] n1102_o;
  wire [8:0] n1104_o;
  wire [8:0] n1105_o;
  wire [8:0] n1107_o;
  wire [8:0] n1108_o;
  wire [8:0] n1109_o;
  wire [8:0] n1110_o;
  wire n1115_o;
  wire [7:0] n1116_o;
  wire n1118_o;
  wire n1120_o;
  wire n1122_o;
  wire n1124_o;
  wire n1125_o;
  wire [15:0] n1128_o;
  wire n1131_o;
  wire n1133_o;
  wire [15:0] n1134_o;
  wire n1136_o;
  wire n1138_o;
  wire [15:0] n1139_o;
  wire [15:0] n1141_o;
  wire [15:0] n1142_o;
  wire [7:0] n1143_o;
  wire [15:0] n1144_o;
  wire [15:0] n1145_o;
  wire n1147_o;
  wire [15:0] n1149_o;
  wire n1151_o;
  wire [7:0] n1152_o;
  wire [15:0] n1154_o;
  wire n1156_o;
  wire [15:0] n1158_o;
  wire n1160_o;
  wire [7:0] n1161_o;
  wire n1163_o;
  wire [12:0] n1164_o;
  wire [7:0] n1165_o;
  wire [7:0] n1166_o;
  wire [7:0] n1167_o;
  wire [7:0] n1169_o;
  wire [7:0] n1170_o;
  wire [7:0] n1171_o;
  wire [7:0] n1172_o;
  wire [7:0] n1173_o;
  wire [7:0] n1174_o;
  reg [7:0] n1175_o;
  wire [7:0] n1176_o;
  wire [7:0] n1177_o;
  wire [7:0] n1178_o;
  wire [7:0] n1180_o;
  wire [7:0] n1181_o;
  wire [7:0] n1182_o;
  wire [7:0] n1183_o;
  wire [7:0] n1184_o;
  wire [7:0] n1185_o;
  reg [7:0] n1186_o;
  wire [15:0] n1187_o;
  wire [15:0] n1191_o;
  reg [15:0] n1192_q;
  wire [15:0] n1194_o;
  wire [7:0] n1195_o;
  wire [7:0] n1197_o;
  wire [7:0] n1198_o;
  wire [7:0] n1200_o;
  wire n1203_o;
  wire n1204_o;
  wire [23:0] n1207_o;
  wire [31:0] n1208_o;
  wire [32:0] n1209_o;
  wire [33:0] n1210_o;
  wire [34:0] n1211_o;
  wire [35:0] n1212_o;
  wire [36:0] n1213_o;
  wire [37:0] n1214_o;
  wire [38:0] n1215_o;
  wire [39:0] n1216_o;
  wire [47:0] n1217_o;
  wire [55:0] n1218_o;
  wire [63:0] n1219_o;
  wire [43:0] n1223_o;
  wire [43:0] n1224_o;
  wire [43:0] n1225_o;
  wire [43:0] n1226_o;
  wire [43:0] n1227_o;
  wire [43:0] n1228_o;
  wire [43:0] n1229_o;
  wire [43:0] n1230_o;
  wire [43:0] n1231_o;
  wire [43:0] n1232_o;
  wire [43:0] n1233_o;
  wire [43:0] n1234_o;
  wire [43:0] n1235_o;
  wire [43:0] n1236_o;
  wire [43:0] n1237_o;
  wire [43:0] n1238_o;
  wire [43:0] n1239_o;
  wire [43:0] n1240_o;
  wire [43:0] n1241_o;
  wire [43:0] n1242_o;
  wire [43:0] n1243_o;
  wire [43:0] n1244_o;
  wire [43:0] n1245_o;
  wire [43:0] n1246_o;
  wire [43:0] n1247_o;
  wire [43:0] n1248_o;
  wire [43:0] n1249_o;
  wire [43:0] n1250_o;
  wire [43:0] n1251_o;
  wire [43:0] n1252_o;
  wire [43:0] n1253_o;
  wire [43:0] n1254_o;
  wire [43:0] n1255_o;
  wire [43:0] n1256_o;
  wire [43:0] n1257_o;
  wire [43:0] n1258_o;
  wire [43:0] n1259_o;
  wire [43:0] n1260_o;
  wire [43:0] n1261_o;
  wire [43:0] n1262_o;
  wire [43:0] n1263_o;
  wire [43:0] n1264_o;
  wire [43:0] n1265_o;
  wire [43:0] n1266_o;
  wire [43:0] n1267_o;
  wire [43:0] n1268_o;
  wire [43:0] n1269_o;
  wire [43:0] n1270_o;
  wire [43:0] n1271_o;
  wire [43:0] n1272_o;
  wire [43:0] n1273_o;
  wire [43:0] n1274_o;
  wire [43:0] n1275_o;
  wire [43:0] n1276_o;
  wire [43:0] n1277_o;
  wire [43:0] n1278_o;
  wire [43:0] n1279_o;
  wire [43:0] n1280_o;
  wire [43:0] n1281_o;
  wire [43:0] n1282_o;
  wire [43:0] n1283_o;
  wire [43:0] n1284_o;
  wire [43:0] n1285_o;
  wire [43:0] n1286_o;
  wire [43:0] n1287_o;
  wire [43:0] n1288_o;
  wire [43:0] n1289_o;
  wire [43:0] n1290_o;
  wire [43:0] n1291_o;
  wire [43:0] n1292_o;
  wire [43:0] n1293_o;
  wire [43:0] n1294_o;
  wire [43:0] n1295_o;
  wire [43:0] n1296_o;
  wire [43:0] n1297_o;
  wire [43:0] n1298_o;
  wire [43:0] n1299_o;
  wire [43:0] n1300_o;
  wire [43:0] n1301_o;
  wire [43:0] n1302_o;
  wire [43:0] n1303_o;
  wire [43:0] n1304_o;
  wire [43:0] n1305_o;
  wire [43:0] n1306_o;
  wire [43:0] n1307_o;
  wire [43:0] n1308_o;
  wire [43:0] n1309_o;
  wire [43:0] n1310_o;
  wire [43:0] n1311_o;
  wire [43:0] n1312_o;
  wire [43:0] n1313_o;
  wire [43:0] n1314_o;
  wire [43:0] n1315_o;
  wire [43:0] n1316_o;
  wire [43:0] n1317_o;
  wire [43:0] n1318_o;
  wire [43:0] n1319_o;
  wire [43:0] n1320_o;
  wire [43:0] n1321_o;
  wire [43:0] n1322_o;
  wire [43:0] n1323_o;
  wire [43:0] n1324_o;
  wire [43:0] n1325_o;
  wire [43:0] n1326_o;
  wire [43:0] n1327_o;
  wire [43:0] n1328_o;
  wire [43:0] n1329_o;
  wire [43:0] n1330_o;
  wire [43:0] n1331_o;
  wire [43:0] n1332_o;
  wire [43:0] n1333_o;
  wire [43:0] n1334_o;
  wire [43:0] n1335_o;
  wire [43:0] n1336_o;
  wire [43:0] n1337_o;
  wire [43:0] n1338_o;
  wire [43:0] n1339_o;
  wire [43:0] n1340_o;
  wire [43:0] n1341_o;
  wire [43:0] n1342_o;
  wire [43:0] n1343_o;
  wire [43:0] n1344_o;
  wire [43:0] n1345_o;
  wire [43:0] n1346_o;
  wire [43:0] n1347_o;
  wire [43:0] n1348_o;
  wire [43:0] n1349_o;
  wire [43:0] n1350_o;
  wire [43:0] n1351_o;
  wire [43:0] n1352_o;
  wire [43:0] n1353_o;
  wire [43:0] n1354_o;
  wire [43:0] n1355_o;
  wire [43:0] n1356_o;
  wire [43:0] n1357_o;
  wire [43:0] n1358_o;
  wire [43:0] n1359_o;
  wire [43:0] n1360_o;
  wire [43:0] n1361_o;
  wire [43:0] n1362_o;
  wire [43:0] n1363_o;
  wire [43:0] n1364_o;
  wire [43:0] n1365_o;
  wire [43:0] n1366_o;
  wire [43:0] n1367_o;
  wire [43:0] n1368_o;
  wire [43:0] n1369_o;
  wire [43:0] n1370_o;
  wire [43:0] n1371_o;
  wire [43:0] n1372_o;
  wire [43:0] n1373_o;
  wire [43:0] n1374_o;
  wire [43:0] n1375_o;
  wire [43:0] n1376_o;
  wire [43:0] n1377_o;
  wire [43:0] n1378_o;
  wire [43:0] n1379_o;
  wire [43:0] n1380_o;
  wire [43:0] n1381_o;
  wire [43:0] n1382_o;
  wire [43:0] n1383_o;
  wire [43:0] n1384_o;
  wire [43:0] n1385_o;
  wire [43:0] n1386_o;
  wire [43:0] n1387_o;
  wire [43:0] n1388_o;
  wire [43:0] n1389_o;
  wire [43:0] n1390_o;
  wire [43:0] n1391_o;
  wire [43:0] n1392_o;
  wire [43:0] n1393_o;
  wire [43:0] n1394_o;
  wire [43:0] n1395_o;
  wire [43:0] n1396_o;
  wire [43:0] n1397_o;
  wire [43:0] n1398_o;
  wire [43:0] n1399_o;
  wire [43:0] n1400_o;
  wire [43:0] n1401_o;
  wire [43:0] n1402_o;
  wire [43:0] n1403_o;
  wire [43:0] n1404_o;
  wire [43:0] n1405_o;
  wire [43:0] n1406_o;
  wire [43:0] n1407_o;
  wire [43:0] n1408_o;
  wire [43:0] n1409_o;
  wire [43:0] n1410_o;
  wire [43:0] n1411_o;
  wire [43:0] n1412_o;
  wire [43:0] n1413_o;
  wire [43:0] n1414_o;
  wire [43:0] n1415_o;
  wire [43:0] n1416_o;
  wire [43:0] n1417_o;
  wire [43:0] n1418_o;
  wire [43:0] n1419_o;
  wire [43:0] n1420_o;
  wire [43:0] n1421_o;
  wire [43:0] n1422_o;
  wire [43:0] n1423_o;
  wire [43:0] n1424_o;
  wire [43:0] n1425_o;
  wire [43:0] n1426_o;
  wire [43:0] n1427_o;
  wire [43:0] n1428_o;
  wire [43:0] n1429_o;
  wire [43:0] n1430_o;
  wire [43:0] n1431_o;
  wire [43:0] n1432_o;
  wire [43:0] n1433_o;
  wire [43:0] n1434_o;
  wire [43:0] n1435_o;
  wire [43:0] n1436_o;
  wire [43:0] n1437_o;
  wire [43:0] n1438_o;
  wire [43:0] n1439_o;
  wire [43:0] n1440_o;
  wire [43:0] n1441_o;
  wire [43:0] n1442_o;
  wire [43:0] n1443_o;
  wire [43:0] n1444_o;
  wire [43:0] n1445_o;
  wire [43:0] n1446_o;
  wire [43:0] n1447_o;
  wire [43:0] n1448_o;
  wire [43:0] n1449_o;
  wire [43:0] n1450_o;
  wire [43:0] n1451_o;
  wire [43:0] n1452_o;
  wire [43:0] n1453_o;
  wire [43:0] n1454_o;
  wire [43:0] n1455_o;
  wire [43:0] n1456_o;
  wire [43:0] n1457_o;
  wire [43:0] n1458_o;
  wire [43:0] n1459_o;
  wire [43:0] n1460_o;
  wire [43:0] n1461_o;
  wire [43:0] n1462_o;
  wire [43:0] n1463_o;
  wire [43:0] n1464_o;
  wire [43:0] n1465_o;
  wire [43:0] n1466_o;
  wire [43:0] n1467_o;
  wire [43:0] n1468_o;
  wire [43:0] n1469_o;
  wire [43:0] n1470_o;
  wire [43:0] n1471_o;
  wire [43:0] n1472_o;
  wire [43:0] n1473_o;
  wire [43:0] n1474_o;
  wire [43:0] n1475_o;
  wire [43:0] n1476_o;
  wire [43:0] n1477_o;
  wire [43:0] n1478_o;
  wire [1:0] n1479_o;
  reg [43:0] n1480_o;
  wire [1:0] n1481_o;
  reg [43:0] n1482_o;
  wire [1:0] n1483_o;
  reg [43:0] n1484_o;
  wire [1:0] n1485_o;
  reg [43:0] n1486_o;
  wire [1:0] n1487_o;
  reg [43:0] n1488_o;
  wire [1:0] n1489_o;
  reg [43:0] n1490_o;
  wire [1:0] n1491_o;
  reg [43:0] n1492_o;
  wire [1:0] n1493_o;
  reg [43:0] n1494_o;
  wire [1:0] n1495_o;
  reg [43:0] n1496_o;
  wire [1:0] n1497_o;
  reg [43:0] n1498_o;
  wire [1:0] n1499_o;
  reg [43:0] n1500_o;
  wire [1:0] n1501_o;
  reg [43:0] n1502_o;
  wire [1:0] n1503_o;
  reg [43:0] n1504_o;
  wire [1:0] n1505_o;
  reg [43:0] n1506_o;
  wire [1:0] n1507_o;
  reg [43:0] n1508_o;
  wire [1:0] n1509_o;
  reg [43:0] n1510_o;
  wire [1:0] n1511_o;
  reg [43:0] n1512_o;
  wire [1:0] n1513_o;
  reg [43:0] n1514_o;
  wire [1:0] n1515_o;
  reg [43:0] n1516_o;
  wire [1:0] n1517_o;
  reg [43:0] n1518_o;
  wire [1:0] n1519_o;
  reg [43:0] n1520_o;
  wire [1:0] n1521_o;
  reg [43:0] n1522_o;
  wire [1:0] n1523_o;
  reg [43:0] n1524_o;
  wire [1:0] n1525_o;
  reg [43:0] n1526_o;
  wire [1:0] n1527_o;
  reg [43:0] n1528_o;
  wire [1:0] n1529_o;
  reg [43:0] n1530_o;
  wire [1:0] n1531_o;
  reg [43:0] n1532_o;
  wire [1:0] n1533_o;
  reg [43:0] n1534_o;
  wire [1:0] n1535_o;
  reg [43:0] n1536_o;
  wire [1:0] n1537_o;
  reg [43:0] n1538_o;
  wire [1:0] n1539_o;
  reg [43:0] n1540_o;
  wire [1:0] n1541_o;
  reg [43:0] n1542_o;
  wire [1:0] n1543_o;
  reg [43:0] n1544_o;
  wire [1:0] n1545_o;
  reg [43:0] n1546_o;
  wire [1:0] n1547_o;
  reg [43:0] n1548_o;
  wire [1:0] n1549_o;
  reg [43:0] n1550_o;
  wire [1:0] n1551_o;
  reg [43:0] n1552_o;
  wire [1:0] n1553_o;
  reg [43:0] n1554_o;
  wire [1:0] n1555_o;
  reg [43:0] n1556_o;
  wire [1:0] n1557_o;
  reg [43:0] n1558_o;
  wire [1:0] n1559_o;
  reg [43:0] n1560_o;
  wire [1:0] n1561_o;
  reg [43:0] n1562_o;
  wire [1:0] n1563_o;
  reg [43:0] n1564_o;
  wire [1:0] n1565_o;
  reg [43:0] n1566_o;
  wire [1:0] n1567_o;
  reg [43:0] n1568_o;
  wire [1:0] n1569_o;
  reg [43:0] n1570_o;
  wire [1:0] n1571_o;
  reg [43:0] n1572_o;
  wire [1:0] n1573_o;
  reg [43:0] n1574_o;
  wire [1:0] n1575_o;
  reg [43:0] n1576_o;
  wire [1:0] n1577_o;
  reg [43:0] n1578_o;
  wire [1:0] n1579_o;
  reg [43:0] n1580_o;
  wire [1:0] n1581_o;
  reg [43:0] n1582_o;
  wire [1:0] n1583_o;
  reg [43:0] n1584_o;
  wire [1:0] n1585_o;
  reg [43:0] n1586_o;
  wire [1:0] n1587_o;
  reg [43:0] n1588_o;
  wire [1:0] n1589_o;
  reg [43:0] n1590_o;
  wire [1:0] n1591_o;
  reg [43:0] n1592_o;
  wire [1:0] n1593_o;
  reg [43:0] n1594_o;
  wire [1:0] n1595_o;
  reg [43:0] n1596_o;
  wire [1:0] n1597_o;
  reg [43:0] n1598_o;
  wire [1:0] n1599_o;
  reg [43:0] n1600_o;
  wire [1:0] n1601_o;
  reg [43:0] n1602_o;
  wire [1:0] n1603_o;
  reg [43:0] n1604_o;
  wire [1:0] n1605_o;
  reg [43:0] n1606_o;
  wire [1:0] n1607_o;
  reg [43:0] n1608_o;
  wire [1:0] n1609_o;
  reg [43:0] n1610_o;
  wire [1:0] n1611_o;
  reg [43:0] n1612_o;
  wire [1:0] n1613_o;
  reg [43:0] n1614_o;
  wire [1:0] n1615_o;
  reg [43:0] n1616_o;
  wire [1:0] n1617_o;
  reg [43:0] n1618_o;
  wire [1:0] n1619_o;
  reg [43:0] n1620_o;
  wire [1:0] n1621_o;
  reg [43:0] n1622_o;
  wire [1:0] n1623_o;
  reg [43:0] n1624_o;
  wire [1:0] n1625_o;
  reg [43:0] n1626_o;
  wire [1:0] n1627_o;
  reg [43:0] n1628_o;
  wire [1:0] n1629_o;
  reg [43:0] n1630_o;
  wire [1:0] n1631_o;
  reg [43:0] n1632_o;
  wire [1:0] n1633_o;
  reg [43:0] n1634_o;
  wire [1:0] n1635_o;
  reg [43:0] n1636_o;
  wire [1:0] n1637_o;
  reg [43:0] n1638_o;
  wire [1:0] n1639_o;
  reg [43:0] n1640_o;
  wire [1:0] n1641_o;
  reg [43:0] n1642_o;
  wire [1:0] n1643_o;
  reg [43:0] n1644_o;
  wire [1:0] n1645_o;
  reg [43:0] n1646_o;
  wire [1:0] n1647_o;
  reg [43:0] n1648_o;
  assign dout= doreg;
  assign addr = myaddr;
  assign nwe = thewe;
  assign sync = n1204_o;
  assign sync_irq = irqactive;
  assign Regs = n1219_o;
  /* R65Cx2.vhd:77:16  */
  assign thecpucycle = n500_q; // (signal)
  /* R65Cx2.vhd:78:16  */
  assign nextcpucycle = n699_o; // (signal)
  /* R65Cx2.vhd:79:16  */
  assign updateregisters = n488_o; // (signal)
  /* R65Cx2.vhd:80:16  */
  assign processirq = n420_q; // (signal)
  /* R65Cx2.vhd:81:16  */
  assign nmireg = n422_q; // (signal)
  /* R65Cx2.vhd:82:16  */
  assign nmiedge = n424_q; // (signal)
  /* R65Cx2.vhd:83:16  */
  assign irqreg = n426_q; // (signal)
  /* R65Cx2.vhd:572:16  */
  assign opcinfo = n453_q; // (signal)
  /* R65Cx2.vhd:573:16  */
  assign nextopcinfo = n1648_o; // (signal)
  /* R65Cx2.vhd:993:134  */
  assign theopcode = n470_q; // (signal)
  /* R65Cx2.vhd:576:16  */
  assign nextopcode = n433_o; // (signal)
  /* R65Cx2.vhd:579:16  */
  assign pc = n973_q; // (signal)
  /* R65Cx2.vhd:598:16  */
  assign nextaddr = n1084_o; // (signal)
  /* R65Cx2.vhd:599:16  */
  assign myaddr = n1192_q; // (signal)
  /* R65Cx2.vhd:600:16  */
  assign myaddrincr = n1194_o; // (signal)
  /* R65Cx2.vhd:601:16  */
  assign myaddrincrh = n1197_o; // (signal)
  /* R65Cx2.vhd:602:16  */
  assign myaddrdecrh = n1200_o; // (signal)
  /* R65Cx2.vhd:603:16  */
  assign thewe = n952_q; // (signal)
  /* R65Cx2.vhd:604:16  */
  assign irqactive = n472_q; // (signal)
  /* R65Cx2.vhd:606:16  */
  assign doreg = n910_q; // (signal)
  /* R65Cx2.vhd:608:16  */
  assign t = n735_q; // (signal)
  /* R65Cx2.vhd:610:16  */
  assign a = n745_q; // (signal)
  /* R65Cx2.vhd:611:16  */
  assign x = n755_q; // (signal)
  /* R65Cx2.vhd:612:16  */
  assign y = n765_q; // (signal)
  /* R65Cx2.vhd:613:16  */
  assign s = n888_q; // (signal)
  /* R65Cx2.vhd:615:16  */
  assign c = n775_q; // (signal)
  /* R65Cx2.vhd:616:16  */
  assign z = n785_q; // (signal)
  /* R65Cx2.vhd:617:16  */
  assign i = n799_q; // (signal)
  /* R65Cx2.vhd:618:16  */
  assign d = n813_q; // (signal)
  /* R65Cx2.vhd:619:16  */
  assign b = 1'bX; // (signal)
  /* R65Cx2.vhd:620:16  */
  assign r = 1'b1; // (signal)
  /* R65Cx2.vhd:621:16  */
  assign v = n823_q; // (signal)
  /* R65Cx2.vhd:622:16  */
  assign n = n833_q; // (signal)
  /* R65Cx2.vhd:735:115  */
  assign aluinput = n32_o; // (signal)
  /* R65Cx2.vhd:627:16  */
  assign alucmpinput = n48_o; // (signal)
  /* R65Cx2.vhd:629:16  */
  assign aluregisterout = n381_o; // (signal)
  /* R65Cx2.vhd:630:16  */
  assign alurmwout = n379_o; // (signal)
  /* R65Cx2.vhd:631:16  */
  assign aluc = n347_o; // (signal)
  /* R65Cx2.vhd:632:16  */
  assign aluz = n377_o; // (signal)
  /* R65Cx2.vhd:633:16  */
  assign aluv = n348_o; // (signal)
  /* R65Cx2.vhd:634:16  */
  assign alun = n378_o; // (signal)
  /* R65Cx2.vhd:636:16  */
  assign indexout = n1110_o; // (signal)
  /* R65Cx2.vhd:645:27  */
  assign n8_o = opcinfo[17];
  /* R65Cx2.vhd:646:38  */
  assign n10_o = 8'b11111111 & a;
  /* R65Cx2.vhd:645:17  */
  assign n12_o = n8_o ? n10_o : 8'b11111111;
  /* R65Cx2.vhd:648:27  */
  assign n14_o = opcinfo[15];
  /* R65Cx2.vhd:649:38  */
  assign n15_o = n12_o & x;
  /* R65Cx2.vhd:648:17  */
  assign n16_o = n14_o ? n15_o : n12_o;
  /* R65Cx2.vhd:651:27  */
  assign n17_o = opcinfo[14];
  /* R65Cx2.vhd:652:38  */
  assign n18_o = n16_o & y;
  /* R65Cx2.vhd:651:17  */
  assign n19_o = n17_o ? n18_o : n16_o;
  /* R65Cx2.vhd:654:27  */
  assign n20_o = opcinfo[13];
  /* R65Cx2.vhd:655:38  */
  assign n21_o = n19_o & s;
  /* R65Cx2.vhd:654:17  */
  assign n22_o = n20_o ? n21_o : n19_o;
  /* R65Cx2.vhd:657:27  */
  assign n23_o = opcinfo[12];
  /* R65Cx2.vhd:658:38  */
  assign n24_o = n22_o & t;
  /* R65Cx2.vhd:657:17  */
  assign n25_o = n23_o ? n24_o : n22_o;
  /* R65Cx2.vhd:660:27  */
  assign n26_o = opcinfo[16];
  /* R65Cx2.vhd:661:38  */
  assign n28_o = n25_o & 8'b11100111;
  /* R65Cx2.vhd:660:17  */
  assign n29_o = n26_o ? n28_o : n25_o;
  /* R65Cx2.vhd:663:27  */
  assign n30_o = opcinfo[10];
  /* R65Cx2.vhd:663:17  */
  assign n32_o = n30_o ? 8'b00000000 : n29_o;
  /* R65Cx2.vhd:675:27  */
  assign n37_o = opcinfo[2];
  /* R65Cx2.vhd:676:38  */
  assign n39_o = 8'b11111111 & a;
  /* R65Cx2.vhd:675:17  */
  assign n41_o = n37_o ? n39_o : 8'b11111111;
  /* R65Cx2.vhd:678:27  */
  assign n43_o = opcinfo[1];
  /* R65Cx2.vhd:679:38  */
  assign n44_o = n41_o & x;
  /* R65Cx2.vhd:678:17  */
  assign n45_o = n43_o ? n44_o : n41_o;
  /* R65Cx2.vhd:681:27  */
  assign n46_o = opcinfo[0];
  /* R65Cx2.vhd:682:38  */
  assign n47_o = n45_o & y;
  /* R65Cx2.vhd:681:17  */
  assign n48_o = n46_o ? n47_o : n45_o;
  /* R65Cx2.vhd:726:29  */
  assign n60_o = opcinfo[9:6];
  /* R65Cx2.vhd:727:70  */
  assign n61_o = {c, aluinput};
  /* R65Cx2.vhd:727:17  */
  assign n63_o = n60_o == 4'b0000;
  /* R65Cx2.vhd:728:78  */
  assign n64_o = {c, n};
  /* R65Cx2.vhd:728:82  */
  assign n65_o = {n64_o, v};
  /* R65Cx2.vhd:728:86  */
  assign n66_o = {n65_o, r};
  /* R65Cx2.vhd:728:93  */
  assign n67_o = ~irqactive;
  /* R65Cx2.vhd:728:90  */
  assign n68_o = {n66_o, n67_o};
  /* R65Cx2.vhd:728:108  */
  assign n69_o = {n68_o, d};
  /* R65Cx2.vhd:728:112  */
  assign n70_o = {n69_o, i};
  /* R65Cx2.vhd:728:116  */
  assign n71_o = {n70_o, z};
  /* R65Cx2.vhd:728:120  */
  assign n72_o = {n71_o, c};
  /* R65Cx2.vhd:728:17  */
  assign n74_o = n60_o == 4'b0001;
  /* R65Cx2.vhd:729:82  */
  assign n76_o = aluinput + 8'b00000001;
  /* R65Cx2.vhd:729:70  */
  assign n77_o = {c, n76_o};
  /* R65Cx2.vhd:729:17  */
  assign n79_o = n60_o == 4'b0010;
  /* R65Cx2.vhd:730:82  */
  assign n81_o = aluinput - 8'b00000001;
  /* R65Cx2.vhd:730:70  */
  assign n82_o = {c, n81_o};
  /* R65Cx2.vhd:730:17  */
  assign n84_o = n60_o == 4'b0011;
  /* R65Cx2.vhd:731:72  */
  assign n86_o = {aluinput, 1'b0};
  /* R65Cx2.vhd:731:17  */
  assign n88_o = n60_o == 4'b1010;
  /* R65Cx2.vhd:732:96  */
  assign n89_o = aluinput | a;
  /* R65Cx2.vhd:732:72  */
  assign n91_o = {1'b0, n89_o};
  /* R65Cx2.vhd:733:128  */
  assign n92_o = aluinput & a;
  /* R65Cx2.vhd:733:104  */
  assign n94_o = {1'b0, n92_o};
  /* R65Cx2.vhd:732:17  */
  assign n96_o = n60_o == 4'b1100;
  /* R65Cx2.vhd:734:96  */
  assign n97_o = ~a;
  /* R65Cx2.vhd:734:91  */
  assign n98_o = aluinput & n97_o;
  /* R65Cx2.vhd:734:67  */
  assign n100_o = {1'b0, n98_o};
  /* R65Cx2.vhd:735:128  */
  assign n101_o = aluinput & a;
  /* R65Cx2.vhd:735:104  */
  assign n103_o = {1'b0, n101_o};
  /* R65Cx2.vhd:734:17  */
  assign n105_o = n60_o == 4'b1101;
  /* R65Cx2.vhd:736:76  */
  assign n106_o = aluinput[0];
  /* R65Cx2.vhd:736:80  */
  assign n107_o = {n106_o, aluinput};
  /* R65Cx2.vhd:736:17  */
  assign n109_o = n60_o == 4'b0100;
  /* R65Cx2.vhd:737:76  */
  assign n110_o = aluinput[0];
  /* R65Cx2.vhd:737:80  */
  assign n112_o = {n110_o, 1'b0};
  /* R65Cx2.vhd:737:96  */
  assign n113_o = aluinput[7:1];
  /* R65Cx2.vhd:737:86  */
  assign n114_o = {n112_o, n113_o};
  /* R65Cx2.vhd:737:17  */
  assign n116_o = n60_o == 4'b1000;
  /* R65Cx2.vhd:738:77  */
  assign n117_o = {aluinput, c};
  /* R65Cx2.vhd:738:17  */
  assign n119_o = n60_o == 4'b1011;
  /* R65Cx2.vhd:739:76  */
  assign n120_o = aluinput[0];
  /* R65Cx2.vhd:739:80  */
  assign n121_o = {n120_o, c};
  /* R65Cx2.vhd:739:94  */
  assign n122_o = aluinput[7:1];
  /* R65Cx2.vhd:739:84  */
  assign n123_o = {n121_o, n122_o};
  /* R65Cx2.vhd:739:17  */
  assign n125_o = n60_o == 4'b1001;
  /* R65Cx2.vhd:740:78  */
  assign n126_o = {c, aluinput};
  assign n127_o = {n125_o, n119_o, n116_o, n109_o, n105_o, n96_o, n88_o, n84_o, n79_o, n74_o, n63_o};
  /* R65Cx2.vhd:726:17  */
  always @*
    case (n127_o)
      11'b10000000000: n128_o <= n123_o;
      11'b01000000000: n128_o <= n117_o;
      11'b00100000000: n128_o <= n114_o;
      11'b00010000000: n128_o <= n107_o;
      11'b00001000000: n128_o <= n100_o;
      11'b00000100000: n128_o <= n91_o;
      11'b00000010000: n128_o <= n86_o;
      11'b00000001000: n128_o <= n82_o;
      11'b00000000100: n128_o <= n77_o;
      11'b00000000010: n128_o <= n72_o;
      11'b00000000001: n128_o <= n61_o;
    endcase
  /* R65Cx2.vhd:726:17  */
  always @*
    case (n127_o)
      11'b10000000000: n131_o <= 9'bXXXXXXXXX;
      11'b01000000000: n131_o <= 9'bXXXXXXXXX;
      11'b00100000000: n131_o <= 9'bXXXXXXXXX;
      11'b00010000000: n131_o <= 9'bXXXXXXXXX;
      11'b00001000000: n131_o <= n103_o;
      11'b00000100000: n131_o <= n94_o;
      11'b00000010000: n131_o <= 9'bXXXXXXXXX;
      11'b00000001000: n131_o <= 9'bXXXXXXXXX;
      11'b00000000100: n131_o <= 9'bXXXXXXXXX;
      11'b00000000010: n131_o <= 9'bXXXXXXXXX;
      11'b00000000001: n131_o <= 9'bXXXXXXXXX;
    endcase
  /* R65Cx2.vhd:744:29  */
  assign n133_o = opcinfo[5:3];
  /* R65Cx2.vhd:745:76  */
  assign n134_o = a[3:0];
  /* R65Cx2.vhd:745:73  */
  assign n136_o = {1'b0, n134_o};
  /* R65Cx2.vhd:745:98  */
  assign n137_o = n128_o[8];
  /* R65Cx2.vhd:745:89  */
  assign n138_o = {n136_o, n137_o};
  /* R65Cx2.vhd:745:119  */
  assign n139_o = n128_o[3:0];
  /* R65Cx2.vhd:745:110  */
  assign n141_o = {1'b0, n139_o};
  /* R65Cx2.vhd:745:132  */
  assign n143_o = {n141_o, 1'b1};
  /* R65Cx2.vhd:745:103  */
  assign n144_o = n138_o + n143_o;
  /* R65Cx2.vhd:746:106  */
  assign n146_o = {1'b0, a};
  /* R65Cx2.vhd:746:127  */
  assign n147_o = n128_o[7:0];
  /* R65Cx2.vhd:746:118  */
  assign n149_o = {1'b0, n147_o};
  /* R65Cx2.vhd:746:111  */
  assign n150_o = n146_o + n149_o;
  /* R65Cx2.vhd:746:165  */
  assign n151_o = n128_o[8];
  /* R65Cx2.vhd:746:156  */
  assign n153_o = {8'b00000000, n151_o};
  /* R65Cx2.vhd:746:141  */
  assign n154_o = n150_o + n153_o;
  /* R65Cx2.vhd:745:17  */
  assign n156_o = n133_o == 3'b010;
  /* R65Cx2.vhd:747:76  */
  assign n157_o = a[3:0];
  /* R65Cx2.vhd:747:73  */
  assign n159_o = {1'b0, n157_o};
  /* R65Cx2.vhd:747:98  */
  assign n160_o = n128_o[8];
  /* R65Cx2.vhd:747:89  */
  assign n161_o = {n159_o, n160_o};
  /* R65Cx2.vhd:747:124  */
  assign n162_o = n128_o[3:0];
  /* R65Cx2.vhd:747:113  */
  assign n163_o = ~n162_o;
  /* R65Cx2.vhd:747:110  */
  assign n165_o = {1'b0, n163_o};
  /* R65Cx2.vhd:747:138  */
  assign n167_o = {n165_o, 1'b1};
  /* R65Cx2.vhd:747:103  */
  assign n168_o = n161_o + n167_o;
  /* R65Cx2.vhd:748:106  */
  assign n170_o = {1'b0, a};
  /* R65Cx2.vhd:748:132  */
  assign n171_o = n128_o[7:0];
  /* R65Cx2.vhd:748:121  */
  assign n172_o = ~n171_o;
  /* R65Cx2.vhd:748:118  */
  assign n174_o = {1'b0, n172_o};
  /* R65Cx2.vhd:748:111  */
  assign n175_o = n170_o + n174_o;
  /* R65Cx2.vhd:748:171  */
  assign n176_o = n128_o[8];
  /* R65Cx2.vhd:748:162  */
  assign n178_o = {8'b00000000, n176_o};
  /* R65Cx2.vhd:748:147  */
  assign n179_o = n175_o + n178_o;
  /* R65Cx2.vhd:747:17  */
  assign n181_o = n133_o == 3'b011;
  /* R65Cx2.vhd:749:74  */
  assign n183_o = {1'b0, alucmpinput};
  /* R65Cx2.vhd:749:110  */
  assign n184_o = n128_o[7:0];
  /* R65Cx2.vhd:749:99  */
  assign n185_o = ~n184_o;
  /* R65Cx2.vhd:749:96  */
  assign n187_o = {1'b0, n185_o};
  /* R65Cx2.vhd:749:89  */
  assign n188_o = n183_o + n187_o;
  /* R65Cx2.vhd:749:125  */
  assign n190_o = n188_o + 9'b000000001;
  /* R65Cx2.vhd:749:17  */
  assign n192_o = n133_o == 3'b001;
  /* R65Cx2.vhd:750:76  */
  assign n193_o = n128_o[8];
  /* R65Cx2.vhd:750:96  */
  assign n194_o = n128_o[7:0];
  /* R65Cx2.vhd:750:85  */
  assign n195_o = a & n194_o;
  /* R65Cx2.vhd:750:80  */
  assign n196_o = {n193_o, n195_o};
  /* R65Cx2.vhd:750:17  */
  assign n198_o = n133_o == 3'b100;
  /* R65Cx2.vhd:751:76  */
  assign n199_o = n128_o[8];
  /* R65Cx2.vhd:751:96  */
  assign n200_o = n128_o[7:0];
  /* R65Cx2.vhd:751:85  */
  assign n201_o = a ^ n200_o;
  /* R65Cx2.vhd:751:80  */
  assign n202_o = {n199_o, n201_o};
  /* R65Cx2.vhd:751:17  */
  assign n204_o = n133_o == 3'b110;
  /* R65Cx2.vhd:752:76  */
  assign n205_o = n128_o[8];
  /* R65Cx2.vhd:752:95  */
  assign n206_o = n128_o[7:0];
  /* R65Cx2.vhd:752:85  */
  assign n207_o = a | n206_o;
  /* R65Cx2.vhd:752:80  */
  assign n208_o = {n205_o, n207_o};
  /* R65Cx2.vhd:752:17  */
  assign n210_o = n133_o == 3'b101;
  /* R65Cx2.vhd:753:17  */
  assign n212_o = n133_o == 3'b111;
  assign n213_o = {n212_o, n210_o, n204_o, n198_o, n192_o, n181_o, n156_o};
  /* R65Cx2.vhd:744:17  */
  always @*
    case (n213_o)
      7'b1000000: n215_o <= 6'bXXXXXX;
      7'b0100000: n215_o <= 6'bXXXXXX;
      7'b0010000: n215_o <= 6'bXXXXXX;
      7'b0001000: n215_o <= 6'bXXXXXX;
      7'b0000100: n215_o <= 6'bXXXXXX;
      7'b0000010: n215_o <= n168_o;
      7'b0000001: n215_o <= n144_o;
    endcase
  /* R65Cx2.vhd:744:17  */
  always @*
    case (n213_o)
      7'b1000000: n218_o <= 9'b000110000;
      7'b0100000: n218_o <= n208_o;
      7'b0010000: n218_o <= n202_o;
      7'b0001000: n218_o <= n196_o;
      7'b0000100: n218_o <= n190_o;
      7'b0000010: n218_o <= n179_o;
      7'b0000001: n218_o <= n154_o;
    endcase
  /* R65Cx2.vhd:758:33  */
  assign n220_o = aluinput[6];
  /* R65Cx2.vhd:761:28  */
  assign n221_o = opcinfo[9:6];
  /* R65Cx2.vhd:761:57  */
  assign n223_o = n221_o == 4'b0100;
  /* R65Cx2.vhd:762:40  */
  assign n224_o = n128_o[1];
  /* R65Cx2.vhd:763:31  */
  assign n225_o = opcinfo[9:6];
  /* R65Cx2.vhd:763:60  */
  assign n227_o = n225_o == 4'b1100;
  /* R65Cx2.vhd:763:85  */
  assign n228_o = opcinfo[9:6];
  /* R65Cx2.vhd:763:114  */
  assign n230_o = n228_o == 4'b1101;
  /* R65Cx2.vhd:763:74  */
  assign n231_o = n227_o | n230_o;
  /* R65Cx2.vhd:764:51  */
  assign n232_o = n131_o[7:0];
  /* R65Cx2.vhd:764:64  */
  assign n234_o = n232_o == 8'b00000000;
  /* R65Cx2.vhd:764:41  */
  assign n237_o = n234_o ? 1'b1 : 1'b0;
  /* R65Cx2.vhd:769:31  */
  assign n238_o = n218_o[7:0];
  /* R65Cx2.vhd:769:44  */
  assign n240_o = n238_o == 8'b00000000;
  /* R65Cx2.vhd:769:17  */
  assign n243_o = n240_o ? 1'b1 : 1'b0;
  /* R65Cx2.vhd:763:17  */
  assign n244_o = n231_o ? n237_o : n243_o;
  /* R65Cx2.vhd:761:17  */
  assign n245_o = n223_o ? n224_o : n244_o;
  /* R65Cx2.vhd:775:28  */
  assign n246_o = opcinfo[9:6];
  /* R65Cx2.vhd:775:57  */
  assign n248_o = n246_o == 4'b0101;
  /* R65Cx2.vhd:775:82  */
  assign n249_o = opcinfo[9:6];
  /* R65Cx2.vhd:775:111  */
  assign n251_o = n249_o == 4'b0100;
  /* R65Cx2.vhd:775:71  */
  assign n252_o = n248_o | n251_o;
  /* R65Cx2.vhd:776:40  */
  assign n253_o = n128_o[7];
  /* R65Cx2.vhd:778:41  */
  assign n254_o = n218_o[7];
  /* R65Cx2.vhd:775:17  */
  assign n255_o = n252_o ? n253_o : n254_o;
  /* R65Cx2.vhd:781:33  */
  assign n256_o = n218_o[8];
  /* R65Cx2.vhd:783:29  */
  assign n257_o = opcinfo[5:3];
  /* R65Cx2.vhd:793:43  */
  assign n258_o = n215_o[5:1];
  /* R65Cx2.vhd:793:56  */
  assign n260_o = $unsigned(n258_o) > $unsigned(5'b01001);
  /* R65Cx2.vhd:794:73  */
  assign n261_o = n218_o[3:0];
  /* R65Cx2.vhd:794:86  */
  assign n263_o = n261_o + 4'b0110;
  /* R65Cx2.vhd:795:51  */
  assign n264_o = n215_o[5];
  /* R65Cx2.vhd:795:55  */
  assign n265_o = ~n264_o;
  assign n266_o = n218_o[8:4];
  assign n267_o = {n266_o, n263_o};
  /* R65Cx2.vhd:796:81  */
  assign n268_o = n267_o[8:4];
  /* R65Cx2.vhd:796:94  */
  assign n270_o = n268_o + 5'b00001;
  assign n271_o = n218_o[8:4];
  /* R65Cx2.vhd:795:41  */
  assign n272_o = n265_o ? n270_o : n271_o;
  assign n273_o = {n272_o, n263_o};
  /* R65Cx2.vhd:792:25  */
  assign n274_o = n275_o ? n273_o : n218_o;
  /* R65Cx2.vhd:792:25  */
  assign n275_o = d & n260_o;
  /* R65Cx2.vhd:790:17  */
  assign n277_o = n257_o == 3'b010;
  /* R65Cx2.vhd:783:17  */
  always @*
    case (n277_o)
      1'b1: n278_o <= n274_o;
    endcase
  /* R65Cx2.vhd:803:29  */
  assign n279_o = opcinfo[5:3];
  /* R65Cx2.vhd:806:35  */
  assign n280_o = a[7];
  /* R65Cx2.vhd:806:51  */
  assign n281_o = n278_o[7];
  /* R65Cx2.vhd:806:39  */
  assign n282_o = n280_o ^ n281_o;
  /* R65Cx2.vhd:806:68  */
  assign n283_o = n128_o[7];
  /* R65Cx2.vhd:806:84  */
  assign n284_o = n278_o[7];
  /* R65Cx2.vhd:806:72  */
  assign n285_o = n283_o ^ n284_o;
  /* R65Cx2.vhd:806:56  */
  assign n286_o = n282_o & n285_o;
  /* R65Cx2.vhd:808:44  */
  assign n287_o = n278_o[8:4];
  /* R65Cx2.vhd:808:57  */
  assign n289_o = $unsigned(n287_o) > $unsigned(5'b01001);
  /* R65Cx2.vhd:809:73  */
  assign n290_o = n278_o[8:4];
  /* R65Cx2.vhd:809:86  */
  assign n292_o = n290_o + 5'b00110;
  assign n293_o = n278_o[8:4];
  /* R65Cx2.vhd:807:25  */
  assign n294_o = n298_o ? n292_o : n293_o;
  /* R65Cx2.vhd:807:25  */
  assign n296_o = n299_o ? 1'b1 : n256_o;
  /* R65Cx2.vhd:807:25  */
  assign n298_o = d & n289_o;
  /* R65Cx2.vhd:807:25  */
  assign n299_o = d & n289_o;
  /* R65Cx2.vhd:804:17  */
  assign n301_o = n279_o == 3'b010;
  /* R65Cx2.vhd:815:35  */
  assign n302_o = a[7];
  /* R65Cx2.vhd:815:51  */
  assign n303_o = n278_o[7];
  /* R65Cx2.vhd:815:39  */
  assign n304_o = n302_o ^ n303_o;
  /* R65Cx2.vhd:815:73  */
  assign n305_o = n128_o[7];
  /* R65Cx2.vhd:815:62  */
  assign n306_o = ~n305_o;
  /* R65Cx2.vhd:815:90  */
  assign n307_o = n278_o[7];
  /* R65Cx2.vhd:815:78  */
  assign n308_o = n306_o ^ n307_o;
  /* R65Cx2.vhd:815:56  */
  assign n309_o = n304_o & n308_o;
  /* R65Cx2.vhd:818:43  */
  assign n310_o = n215_o[5];
  /* R65Cx2.vhd:818:47  */
  assign n311_o = ~n310_o;
  /* R65Cx2.vhd:819:73  */
  assign n312_o = n278_o[7:0];
  /* R65Cx2.vhd:819:86  */
  assign n314_o = n312_o - 8'b00000110;
  assign n315_o = n278_o[7:0];
  /* R65Cx2.vhd:818:33  */
  assign n316_o = n311_o ? n314_o : n315_o;
  assign n317_o = n278_o[8];
  assign n318_o = {n317_o, n316_o};
  /* R65Cx2.vhd:822:44  */
  assign n319_o = n318_o[8];
  /* R65Cx2.vhd:822:48  */
  assign n320_o = ~n319_o;
  assign n321_o = n278_o[8];
  assign n322_o = {n321_o, n316_o};
  /* R65Cx2.vhd:823:73  */
  assign n323_o = n322_o[8:4];
  /* R65Cx2.vhd:823:86  */
  assign n325_o = n323_o - 5'b00110;
  assign n326_o = n314_o[7:4];
  assign n327_o = n278_o[7:4];
  /* R65Cx2.vhd:818:33  */
  assign n328_o = n311_o ? n326_o : n327_o;
  assign n329_o = n278_o[8];
  assign n330_o = {n329_o, n328_o};
  /* R65Cx2.vhd:822:33  */
  assign n331_o = n320_o ? n325_o : n330_o;
  assign n332_o = n314_o[3:0];
  assign n333_o = n278_o[3:0];
  /* R65Cx2.vhd:818:33  */
  assign n334_o = n311_o ? n332_o : n333_o;
  assign n335_o = {n331_o, n334_o};
  /* R65Cx2.vhd:816:25  */
  assign n336_o = d ? n335_o : n278_o;
  /* R65Cx2.vhd:814:17  */
  assign n338_o = n279_o == 3'b011;
  assign n339_o = {n338_o, n301_o};
  assign n340_o = n336_o[3:0];
  assign n341_o = n278_o[3:0];
  /* R65Cx2.vhd:803:17  */
  always @*
    case (n339_o)
      2'b10: n342_o <= n340_o;
      2'b01: n342_o <= n341_o;
    endcase
  assign n343_o = n336_o[8:4];
  assign n344_o = n278_o[8:4];
  /* R65Cx2.vhd:803:17  */
  always @*
    case (n339_o)
      2'b10: n345_o <= n343_o;
      2'b01: n345_o <= n294_o;
    endcase
  /* R65Cx2.vhd:803:17  */
  always @*
    case (n339_o)
      2'b10: n347_o <= n256_o;
      2'b01: n347_o <= n296_o;
    endcase
  /* R65Cx2.vhd:803:17  */
  always @*
    case (n339_o)
      2'b10: n348_o <= n309_o;
      2'b01: n348_o <= n286_o;
    endcase
  /* R65Cx2.vhd:830:29  */
  assign n349_o = opcinfo[5:3];
  assign n350_o = {n345_o, n342_o};
  /* R65Cx2.vhd:833:44  */
  assign n351_o = n350_o[7:0];
  /* R65Cx2.vhd:833:57  */
  assign n353_o = n351_o == 8'b00000000;
  /* R65Cx2.vhd:833:33  */
  assign n356_o = n353_o ? 1'b1 : 1'b0;
  assign n357_o = {n345_o, n342_o};
  /* R65Cx2.vhd:838:33  */
  assign n358_o = n357_o[7];
  /* R65Cx2.vhd:832:25  */
  assign n359_o = d ? n356_o : n245_o;
  /* R65Cx2.vhd:832:25  */
  assign n360_o = d ? n358_o : n255_o;
  /* R65Cx2.vhd:831:17  */
  assign n362_o = n349_o == 3'b010;
  assign n363_o = {n345_o, n342_o};
  /* R65Cx2.vhd:842:44  */
  assign n364_o = n363_o[7:0];
  /* R65Cx2.vhd:842:57  */
  assign n366_o = n364_o == 8'b00000000;
  /* R65Cx2.vhd:842:33  */
  assign n369_o = n366_o ? 1'b1 : 1'b0;
  assign n370_o = {n345_o, n342_o};
  /* R65Cx2.vhd:847:33  */
  assign n371_o = n370_o[7];
  /* R65Cx2.vhd:841:25  */
  assign n372_o = d ? n369_o : n245_o;
  /* R65Cx2.vhd:841:25  */
  assign n373_o = d ? n371_o : n255_o;
  /* R65Cx2.vhd:840:17  */
  assign n375_o = n349_o == 3'b011;
  assign n376_o = {n375_o, n362_o};
  /* R65Cx2.vhd:830:17  */
  always @*
    case (n376_o)
      2'b10: n377_o <= n372_o;
      2'b01: n377_o <= n359_o;
    endcase
  /* R65Cx2.vhd:830:17  */
  always @*
    case (n376_o)
      2'b10: n378_o <= n373_o;
      2'b01: n378_o <= n360_o;
    endcase
  /* R65Cx2.vhd:854:37  */
  assign n379_o = n128_o[7:0];
  assign n380_o = {n345_o, n342_o};
  /* R65Cx2.vhd:855:43  */
  assign n381_o = n380_o[7:0];
  /* R65Cx2.vhd:868:48  */
  assign n388_o = thecpucycle == 5'b10000;
  /* R65Cx2.vhd:868:71  */
  assign n389_o = ~reset;
  /* R65Cx2.vhd:868:62  */
  assign n390_o = n388_o | n389_o;
  /* R65Cx2.vhd:868:33  */
  assign n392_o = n390_o ? 1'b1 : nmireg;
  /* R65Cx2.vhd:871:49  */
  assign n394_o = nextcpucycle != 5'b00101;
  /* R65Cx2.vhd:871:90  */
  assign n396_o = nextcpucycle != 5'b00000;
  /* R65Cx2.vhd:871:73  */
  assign n397_o = n394_o & n396_o;
  /* R65Cx2.vhd:874:71  */
  assign n398_o = ~nmi_n;
  /* R65Cx2.vhd:874:60  */
  assign n399_o = nmiedge & n398_o;
  /* R65Cx2.vhd:871:33  */
  assign n401_o = n402_o ? 1'b0 : n392_o;
  /* R65Cx2.vhd:871:33  */
  assign n402_o = n397_o & n399_o;
  /* R65Cx2.vhd:880:72  */
  assign n405_o = irqreg | i;
  /* R65Cx2.vhd:880:60  */
  assign n406_o = nmireg & n405_o;
  /* R65Cx2.vhd:880:89  */
  assign n407_o = opcinfo[18];
  /* R65Cx2.vhd:880:79  */
  assign n408_o = n406_o | n407_o;
  /* R65Cx2.vhd:880:47  */
  assign n409_o = ~n408_o;
  /* R65Cx2.vhd:867:25  */
  assign n412_o = enable & n397_o;
  /* R65Cx2.vhd:867:25  */
  assign n413_o = enable & n397_o;
  /* R65Cx2.vhd:866:17  */
  assign n419_o = enable ? n409_o : processirq;
  /* R65Cx2.vhd:866:17  */
  always @(posedge clk)
    n420_q <= n419_o;
  /* R65Cx2.vhd:866:17  */
  assign n421_o = enable ? n401_o : nmireg;
  /* R65Cx2.vhd:866:17  */
  always @(posedge clk)
    n422_q <= n421_o;
  /* R65Cx2.vhd:866:17  */
  assign n423_o = n412_o ? nmi_n : nmiedge;
  /* R65Cx2.vhd:866:17  */
  always @(posedge clk)
    n424_q <= n423_o;
  /* R65Cx2.vhd:866:17  */
  assign n425_o = n413_o ? irq_n : irqreg;
  /* R65Cx2.vhd:866:17  */
  always @(posedge clk)
    n426_q <= n425_o;
  /* R65Cx2.vhd:904:26  */
  assign n429_o = ~reset;
  /* R65Cx2.vhd:906:17  */
  assign n431_o = processirq ? 8'b00000000 : di;
  /* R65Cx2.vhd:904:17  */
  assign n433_o = n429_o ? 8'b01001100 : n431_o;
  /* R65Cx2.vhd:912:39  */
  assign n438_o = 8'b11111111 - nextopcode;
  /* R65Cx2.vhd:928:43  */
  assign n444_o = ~reset;
  /* R65Cx2.vhd:928:66  */
  assign n446_o = thecpucycle == 5'b00000;
  /* R65Cx2.vhd:928:50  */
  assign n447_o = n444_o | n446_o;
  /* R65Cx2.vhd:927:25  */
  assign n449_o = enable & n447_o;
  /* R65Cx2.vhd:926:17  */
  assign n452_o = n449_o ? nextopcinfo : opcinfo;
  /* R65Cx2.vhd:926:17  */
  always @(posedge clk)
    n453_q <= n452_o;
  /* R65Cx2.vhd:939:48  */
  assign n457_o = thecpucycle == 5'b00000;
  /* R65Cx2.vhd:941:41  */
  assign n460_o = processirq ? 1'b1 : 1'b0;
  /* R65Cx2.vhd:938:25  */
  assign n464_o = enable & n457_o;
  /* R65Cx2.vhd:938:25  */
  assign n465_o = enable & n457_o;
  /* R65Cx2.vhd:937:17  */
  assign n469_o = n464_o ? nextopcode : theopcode;
  /* R65Cx2.vhd:937:17  */
  always @(posedge clk)
    n470_q <= n469_o;
  /* R65Cx2.vhd:937:17  */
  assign n471_o = n465_o ? n460_o : irqactive;
  /* R65Cx2.vhd:937:17  */
  always @(posedge clk)
    n472_q <= n471_o;
  /* R65Cx2.vhd:958:35  */
  assign n475_o = opcinfo[19];
  /* R65Cx2.vhd:959:48  */
  assign n477_o = thecpucycle == 5'b01000;
  /* R65Cx2.vhd:959:33  */
  assign n480_o = n477_o ? 1'b1 : 1'b0;
  /* R65Cx2.vhd:962:43  */
  assign n482_o = thecpucycle == 5'b00000;
  /* R65Cx2.vhd:962:25  */
  assign n485_o = n482_o ? 1'b1 : 1'b0;
  /* R65Cx2.vhd:958:25  */
  assign n486_o = n475_o ? n480_o : n485_o;
  /* R65Cx2.vhd:957:17  */
  assign n488_o = enable ? n486_o : 1'b0;
  /* R65Cx2.vhd:971:25  */
  assign n494_o = enable ? nextcpucycle : thecpucycle;
  /* R65Cx2.vhd:974:34  */
  assign n495_o = ~reset;
  /* R65Cx2.vhd:974:25  */
  assign n497_o = n495_o ? 5'b00001 : n494_o;
  /* R65Cx2.vhd:970:17  */
  always @(posedge clk)
    n500_q <= n497_o;
  /* R65Cx2.vhd:987:17  */
  assign n503_o = thecpucycle == 5'b00000;
  /* R65Cx2.vhd:988:91  */
  assign n504_o = opcinfo[26];
  /* R65Cx2.vhd:989:130  */
  assign n505_o = theopcode[5];
  /* R65Cx2.vhd:989:119  */
  assign n506_o = n == n505_o;
  /* R65Cx2.vhd:989:147  */
  assign n507_o = theopcode[7:6];
  /* R65Cx2.vhd:989:160  */
  assign n509_o = n507_o == 2'b00;
  /* R65Cx2.vhd:989:134  */
  assign n510_o = n506_o & n509_o;
  /* R65Cx2.vhd:990:138  */
  assign n511_o = theopcode[5];
  /* R65Cx2.vhd:990:127  */
  assign n512_o = v == n511_o;
  /* R65Cx2.vhd:990:155  */
  assign n513_o = theopcode[7:6];
  /* R65Cx2.vhd:990:168  */
  assign n515_o = n513_o == 2'b01;
  /* R65Cx2.vhd:990:142  */
  assign n516_o = n512_o & n515_o;
  /* R65Cx2.vhd:990:121  */
  assign n517_o = n510_o | n516_o;
  /* R65Cx2.vhd:991:138  */
  assign n518_o = theopcode[5];
  /* R65Cx2.vhd:991:127  */
  assign n519_o = c == n518_o;
  /* R65Cx2.vhd:991:155  */
  assign n520_o = theopcode[7:6];
  /* R65Cx2.vhd:991:168  */
  assign n522_o = n520_o == 2'b10;
  /* R65Cx2.vhd:991:142  */
  assign n523_o = n519_o & n522_o;
  /* R65Cx2.vhd:991:121  */
  assign n524_o = n517_o | n523_o;
  /* R65Cx2.vhd:992:138  */
  assign n525_o = theopcode[5];
  /* R65Cx2.vhd:992:127  */
  assign n526_o = z == n525_o;
  /* R65Cx2.vhd:992:155  */
  assign n527_o = theopcode[7:6];
  /* R65Cx2.vhd:992:168  */
  assign n529_o = n527_o == 2'b11;
  /* R65Cx2.vhd:992:142  */
  assign n530_o = n526_o & n529_o;
  /* R65Cx2.vhd:992:121  */
  assign n531_o = n524_o | n530_o;
  /* R65Cx2.vhd:993:147  */
  assign n533_o = theopcode == 8'b10000000;
  /* R65Cx2.vhd:993:121  */
  assign n534_o = n531_o | n533_o;
  /* R65Cx2.vhd:989:113  */
  assign n537_o = n534_o ? 5'b00101 : 5'b00000;
  /* R65Cx2.vhd:996:119  */
  assign n538_o = opcinfo[23];
  /* R65Cx2.vhd:998:118  */
  assign n539_o = opcinfo[29];
  /* R65Cx2.vhd:998:156  */
  assign n540_o = opcinfo[28];
  /* R65Cx2.vhd:998:145  */
  assign n541_o = n539_o & n540_o;
  /* R65Cx2.vhd:1000:118  */
  assign n542_o = opcinfo[29];
  /* R65Cx2.vhd:1002:118  */
  assign n543_o = opcinfo[28];
  /* R65Cx2.vhd:1004:118  */
  assign n544_o = opcinfo[32];
  /* R65Cx2.vhd:1006:118  */
  assign n545_o = opcinfo[30];
  /* R65Cx2.vhd:1007:131  */
  assign n546_o = opcinfo[25];
  /* R65Cx2.vhd:1007:121  */
  assign n549_o = n546_o ? 5'b00011 : 5'b00100;
  /* R65Cx2.vhd:1012:118  */
  assign n550_o = opcinfo[31];
  /* R65Cx2.vhd:1013:131  */
  assign n551_o = opcinfo[22];
  /* R65Cx2.vhd:1014:148  */
  assign n552_o = opcinfo[25];
  /* R65Cx2.vhd:1014:180  */
  assign n553_o = opcinfo[24];
  /* R65Cx2.vhd:1014:169  */
  assign n554_o = n552_o | n553_o;
  /* R65Cx2.vhd:1014:137  */
  assign n557_o = n554_o ? 5'b01011 : 5'b01100;
  /* R65Cx2.vhd:1020:148  */
  assign n558_o = opcinfo[25];
  /* R65Cx2.vhd:1020:180  */
  assign n559_o = opcinfo[24];
  /* R65Cx2.vhd:1020:169  */
  assign n560_o = n558_o | n559_o;
  /* R65Cx2.vhd:1020:137  */
  assign n563_o = n560_o ? 5'b00111 : 5'b01001;
  /* R65Cx2.vhd:1013:121  */
  assign n564_o = n551_o ? n557_o : n563_o;
  /* R65Cx2.vhd:1026:118  */
  assign n565_o = opcinfo[27];
  /* R65Cx2.vhd:1026:105  */
  assign n568_o = n565_o ? 5'b10001 : 5'b00000;
  /* R65Cx2.vhd:1012:105  */
  assign n569_o = n550_o ? n564_o : n568_o;
  /* R65Cx2.vhd:1006:105  */
  assign n570_o = n545_o ? n549_o : n569_o;
  /* R65Cx2.vhd:1004:105  */
  assign n572_o = n544_o ? 5'b00010 : n570_o;
  /* R65Cx2.vhd:1002:105  */
  assign n574_o = n543_o ? 5'b01100 : n572_o;
  /* R65Cx2.vhd:1000:105  */
  assign n576_o = n542_o ? 5'b01101 : n574_o;
  /* R65Cx2.vhd:998:105  */
  assign n578_o = n541_o ? 5'b01110 : n576_o;
  /* R65Cx2.vhd:996:105  */
  assign n580_o = n538_o ? 5'b01101 : n578_o;
  /* R65Cx2.vhd:988:81  */
  assign n581_o = n504_o ? n537_o : n580_o;
  /* R65Cx2.vhd:988:17  */
  assign n583_o = thecpucycle == 5'b00001;
  /* R65Cx2.vhd:1030:123  */
  assign n584_o = opcinfo[22];
  /* R65Cx2.vhd:1031:140  */
  assign n585_o = opcinfo[25];
  /* R65Cx2.vhd:1031:172  */
  assign n586_o = opcinfo[24];
  /* R65Cx2.vhd:1031:161  */
  assign n587_o = n585_o | n586_o;
  /* R65Cx2.vhd:1031:129  */
  assign n590_o = n587_o ? 5'b01011 : 5'b01100;
  /* R65Cx2.vhd:1030:113  */
  assign n592_o = n584_o ? n590_o : 5'b01000;
  /* R65Cx2.vhd:1037:124  */
  assign n594_o = opcinfo[30];
  /* R65Cx2.vhd:1037:165  */
  assign n595_o = opcinfo[25];
  /* R65Cx2.vhd:1037:153  */
  assign n596_o = n594_o & n595_o;
  /* R65Cx2.vhd:1038:147  */
  assign n597_o = opcinfo[22];
  /* R65Cx2.vhd:1038:137  */
  assign n600_o = n597_o ? 5'b01100 : 5'b01001;
  /* R65Cx2.vhd:1037:113  */
  assign n601_o = n596_o ? n600_o : n592_o;
  /* R65Cx2.vhd:1029:17  */
  assign n603_o = thecpucycle == 5'b00010;
  /* R65Cx2.vhd:1044:17  */
  assign n605_o = thecpucycle == 5'b00011;
  /* R65Cx2.vhd:1045:17  */
  assign n607_o = thecpucycle == 5'b00100;
  /* R65Cx2.vhd:1046:68  */
  assign n608_o = indexout[8];
  /* R65Cx2.vhd:1046:76  */
  assign n609_o = t[7];
  /* R65Cx2.vhd:1046:72  */
  assign n610_o = n608_o != n609_o;
  /* R65Cx2.vhd:1046:57  */
  assign n613_o = n610_o ? 5'b00110 : 5'b00000;
  /* R65Cx2.vhd:1046:17  */
  assign n615_o = thecpucycle == 5'b00101;
  /* R65Cx2.vhd:1049:75  */
  assign n616_o = opcinfo[31];
  /* R65Cx2.vhd:1049:65  */
  assign n619_o = n616_o ? 5'b01001 : 5'b00000;
  /* R65Cx2.vhd:1049:17  */
  assign n621_o = thecpucycle == 5'b00111;
  /* R65Cx2.vhd:1053:107  */
  assign n622_o = opcinfo[27];
  /* R65Cx2.vhd:1055:111  */
  assign n623_o = indexout[8];
  /* R65Cx2.vhd:1057:110  */
  assign n624_o = opcinfo[21];
  /* R65Cx2.vhd:1059:123  */
  assign n625_o = opcinfo[25];
  /* R65Cx2.vhd:1059:148  */
  assign n626_o = opcinfo[24];
  /* R65Cx2.vhd:1059:138  */
  assign n627_o = n625_o | n626_o;
  /* R65Cx2.vhd:1059:113  */
  assign n630_o = n627_o ? 5'b01001 : 5'b01010;
  /* R65Cx2.vhd:1057:97  */
  assign n633_o = n624_o ? n630_o : 5'b00000;
  /* R65Cx2.vhd:1055:97  */
  assign n635_o = n623_o ? 5'b01001 : n633_o;
  /* R65Cx2.vhd:1053:97  */
  assign n637_o = n622_o ? 5'b10001 : n635_o;
  /* R65Cx2.vhd:1052:17  */
  assign n639_o = thecpucycle == 5'b01000;
  /* R65Cx2.vhd:1063:67  */
  assign n640_o = opcinfo[21];
  /* R65Cx2.vhd:1063:57  */
  assign n643_o = n640_o ? 5'b01010 : 5'b00000;
  /* R65Cx2.vhd:1063:17  */
  assign n645_o = thecpucycle == 5'b01001;
  /* R65Cx2.vhd:1066:17  */
  assign n647_o = thecpucycle == 5'b01010;
  /* R65Cx2.vhd:1067:17  */
  assign n649_o = thecpucycle == 5'b01011;
  /* R65Cx2.vhd:1069:99  */
  assign n650_o = opcinfo[29];
  /* R65Cx2.vhd:1069:89  */
  assign n653_o = n650_o ? 5'b01110 : 5'b01000;
  /* R65Cx2.vhd:1068:17  */
  assign n656_o = thecpucycle == 5'b01101;
  /* R65Cx2.vhd:1073:99  */
  assign n657_o = opcinfo[19];
  /* R65Cx2.vhd:1073:89  */
  assign n660_o = n657_o ? 5'b01000 : 5'b01111;
  /* R65Cx2.vhd:1076:99  */
  assign n662_o = opcinfo[28];
  /* R65Cx2.vhd:1076:114  */
  assign n663_o = ~n662_o;
  /* R65Cx2.vhd:1076:131  */
  assign n664_o = opcinfo[23];
  /* R65Cx2.vhd:1076:120  */
  assign n665_o = n663_o & n664_o;
  /* R65Cx2.vhd:1076:89  */
  assign n667_o = n665_o ? 5'b10001 : n660_o;
  /* R65Cx2.vhd:1072:17  */
  assign n669_o = thecpucycle == 5'b01110;
  /* R65Cx2.vhd:1080:99  */
  assign n670_o = opcinfo[28];
  /* R65Cx2.vhd:1080:114  */
  assign n671_o = ~n670_o;
  /* R65Cx2.vhd:1080:130  */
  assign n672_o = opcinfo[23];
  /* R65Cx2.vhd:1080:120  */
  assign n673_o = n671_o | n672_o;
  /* R65Cx2.vhd:1082:102  */
  assign n674_o = opcinfo[29];
  /* R65Cx2.vhd:1082:89  */
  assign n677_o = n674_o ? 5'b10000 : 5'b01000;
  /* R65Cx2.vhd:1080:89  */
  assign n679_o = n673_o ? 5'b10001 : n677_o;
  /* R65Cx2.vhd:1079:17  */
  assign n682_o = thecpucycle == 5'b01111;
  /* R65Cx2.vhd:1085:17  */
  assign n684_o = thecpucycle == 5'b10000;
  /* R65Cx2.vhd:1086:75  */
  assign n685_o = opcinfo[20];
  /* R65Cx2.vhd:1086:65  */
  assign n688_o = n685_o ? 5'b10010 : 5'b00000;
  /* R65Cx2.vhd:1086:17  */
  assign n690_o = thecpucycle == 5'b10001;
  assign n691_o = {n690_o, n684_o, n682_o, n669_o, n656_o, n649_o, n647_o, n645_o, n639_o, n621_o, n615_o, n607_o, n605_o, n603_o, n583_o, n503_o};
  /* R65Cx2.vhd:986:17  */
  always @*
    case (n691_o)
      16'b1000000000000000: n699_o <= n688_o;
      16'b0100000000000000: n699_o <= 5'b01000;
      16'b0010000000000000: n699_o <= n679_o;
      16'b0001000000000000: n699_o <= n667_o;
      16'b0000100000000000: n699_o <= n653_o;
      16'b0000010000000000: n699_o <= 5'b01100;
      16'b0000001000000000: n699_o <= 5'b01100;
      16'b0000000100000000: n699_o <= n643_o;
      16'b0000000010000000: n699_o <= n637_o;
      16'b0000000001000000: n699_o <= n619_o;
      16'b0000000000100000: n699_o <= n613_o;
      16'b0000000000010000: n699_o <= 5'b00010;
      16'b0000000000001000: n699_o <= 5'b00100;
      16'b0000000000000100: n699_o <= n601_o;
      16'b0000000000000010: n699_o <= n581_o;
      16'b0000000000000001: n699_o <= 5'b00001;
    endcase
  /* R65Cx2.vhd:1101:33  */
  assign n705_o = thecpucycle == 5'b00001;
  /* R65Cx2.vhd:1103:51  */
  assign n706_o = opcinfo[23];
  /* R65Cx2.vhd:1104:70  */
  assign n708_o = theopcode == 8'b00101000;
  /* R65Cx2.vhd:1104:91  */
  assign n710_o = theopcode == 8'b01000000;
  /* R65Cx2.vhd:1104:78  */
  assign n711_o = n708_o | n710_o;
  /* R65Cx2.vhd:1105:74  */
  assign n713_o = di | 8'b00110000;
  /* R65Cx2.vhd:1104:57  */
  assign n714_o = n711_o ? n713_o : di;
  /* R65Cx2.vhd:1103:41  */
  assign n715_o = n706_o ? n714_o : t;
  /* R65Cx2.vhd:1102:33  */
  assign n717_o = thecpucycle == 5'b01101;
  /* R65Cx2.vhd:1102:50  */
  assign n719_o = thecpucycle == 5'b01110;
  /* R65Cx2.vhd:1102:50  */
  assign n720_o = n717_o | n719_o;
  /* R65Cx2.vhd:1110:33  */
  assign n722_o = thecpucycle == 5'b00100;
  /* R65Cx2.vhd:1110:52  */
  assign n724_o = thecpucycle == 5'b01000;
  /* R65Cx2.vhd:1110:52  */
  assign n725_o = n722_o | n724_o;
  /* R65Cx2.vhd:1110:64  */
  assign n727_o = thecpucycle == 5'b01001;
  /* R65Cx2.vhd:1110:64  */
  assign n728_o = n725_o | n727_o;
  assign n729_o = {n728_o, n720_o, n705_o};
  /* R65Cx2.vhd:1100:33  */
  always @*
    case (n729_o)
      3'b100: n730_o <= di;
      3'b010: n730_o <= n715_o;
      3'b001: n730_o <= di;
    endcase
  /* R65Cx2.vhd:1098:17  */
  assign n734_o = enable ? n730_o : t;
  /* R65Cx2.vhd:1098:17  */
  always @(posedge clk)
    n735_q <= n734_o;
  /* R65Cx2.vhd:1124:43  */
  assign n739_o = opcinfo[43];
  /* R65Cx2.vhd:1123:25  */
  assign n741_o = updateregisters & n739_o;
  /* R65Cx2.vhd:1122:17  */
  assign n744_o = n741_o ? aluregisterout : a;
  /* R65Cx2.vhd:1122:17  */
  always @(posedge clk)
    n745_q <= n744_o;
  /* R65Cx2.vhd:1138:43  */
  assign n749_o = opcinfo[42];
  /* R65Cx2.vhd:1137:25  */
  assign n751_o = updateregisters & n749_o;
  /* R65Cx2.vhd:1136:17  */
  assign n754_o = n751_o ? aluregisterout : x;
  /* R65Cx2.vhd:1136:17  */
  always @(posedge clk)
    n755_q <= n754_o;
  /* R65Cx2.vhd:1152:43  */
  assign n759_o = opcinfo[41];
  /* R65Cx2.vhd:1151:25  */
  assign n761_o = updateregisters & n759_o;
  /* R65Cx2.vhd:1150:17  */
  assign n764_o = n761_o ? aluregisterout : y;
  /* R65Cx2.vhd:1150:17  */
  always @(posedge clk)
    n765_q <= n764_o;
  /* R65Cx2.vhd:1166:43  */
  assign n769_o = opcinfo[34];
  /* R65Cx2.vhd:1165:25  */
  assign n771_o = updateregisters & n769_o;
  /* R65Cx2.vhd:1164:17  */
  assign n774_o = n771_o ? aluc : c;
  /* R65Cx2.vhd:1164:17  */
  always @(posedge clk)
    n775_q <= n774_o;
  /* R65Cx2.vhd:1180:43  */
  assign n779_o = opcinfo[35];
  /* R65Cx2.vhd:1179:25  */
  assign n781_o = updateregisters & n779_o;
  /* R65Cx2.vhd:1178:17  */
  assign n784_o = n781_o ? aluz : z;
  /* R65Cx2.vhd:1178:17  */
  always @(posedge clk)
    n785_q <= n784_o;
  /* R65Cx2.vhd:1192:18  */
  assign n788_o = ~reset;
  /* R65Cx2.vhd:1196:43  */
  assign n790_o = opcinfo[36];
  /* R65Cx2.vhd:1197:62  */
  assign n791_o = aluinput[2];
  /* R65Cx2.vhd:1195:25  */
  assign n793_o = updateregisters & n790_o;
  /* R65Cx2.vhd:1194:9  */
  assign n798_o = n793_o ? n791_o : i;
  /* R65Cx2.vhd:1194:9  */
  always @(posedge clk or posedge n788_o)
    if (n788_o)
      n799_q <= 1'b1;
    else
      n799_q <= n798_o;
  /* R65Cx2.vhd:1207:18  */
  assign n802_o = ~reset;
  /* R65Cx2.vhd:1211:43  */
  assign n804_o = opcinfo[37];
  /* R65Cx2.vhd:1212:62  */
  assign n805_o = aluinput[3];
  /* R65Cx2.vhd:1210:25  */
  assign n807_o = updateregisters & n804_o;
  /* R65Cx2.vhd:1209:9  */
  assign n812_o = n807_o ? n805_o : d;
  /* R65Cx2.vhd:1209:9  */
  always @(posedge clk or posedge n802_o)
    if (n802_o)
      n813_q <= 1'b0;
    else
      n813_q <= n812_o;
  /* R65Cx2.vhd:1225:43  */
  assign n817_o = opcinfo[38];
  /* R65Cx2.vhd:1224:25  */
  assign n819_o = updateregisters & n817_o;
  /* R65Cx2.vhd:1223:17  */
  assign n822_o = n819_o ? aluv : v;
  /* R65Cx2.vhd:1223:17  */
  always @(posedge clk)
    n823_q <= n822_o;
  /* R65Cx2.vhd:1239:43  */
  assign n827_o = opcinfo[39];
  /* R65Cx2.vhd:1238:25  */
  assign n829_o = updateregisters & n827_o;
  /* R65Cx2.vhd:1237:17  */
  assign n832_o = n829_o ? alun : n;
  /* R65Cx2.vhd:1237:17  */
  always @(posedge clk)
    n833_q <= n832_o;
  /* R65Cx2.vhd:1255:35  */
  assign n839_o = opcinfo[23];
  /* R65Cx2.vhd:1256:46  */
  assign n841_o = s + 8'b00000001;
  /* R65Cx2.vhd:1258:46  */
  assign n843_o = s - 8'b00000001;
  /* R65Cx2.vhd:1255:25  */
  assign n844_o = n839_o ? n841_o : n843_o;
  /* R65Cx2.vhd:1265:108  */
  assign n845_o = opcinfo[23];
  /* R65Cx2.vhd:1265:139  */
  assign n846_o = opcinfo[28];
  /* R65Cx2.vhd:1265:128  */
  assign n847_o = n845_o | n846_o;
  /* R65Cx2.vhd:1265:97  */
  assign n850_o = n847_o ? 1'b1 : 1'b0;
  /* R65Cx2.vhd:1264:33  */
  assign n852_o = nextcpucycle == 5'b01101;
  /* R65Cx2.vhd:1269:33  */
  assign n854_o = nextcpucycle == 5'b01110;
  /* R65Cx2.vhd:1270:33  */
  assign n856_o = nextcpucycle == 5'b01111;
  /* R65Cx2.vhd:1271:33  */
  assign n858_o = nextcpucycle == 5'b10000;
  /* R65Cx2.vhd:1272:83  */
  assign n859_o = opcinfo[19];
  /* R65Cx2.vhd:1272:73  */
  assign n862_o = n859_o ? 1'b1 : 1'b0;
  /* R65Cx2.vhd:1272:33  */
  assign n864_o = nextcpucycle == 5'b01000;
  /* R65Cx2.vhd:1275:75  */
  assign n865_o = opcinfo[28];
  /* R65Cx2.vhd:1275:65  */
  assign n868_o = n865_o ? 1'b1 : 1'b0;
  /* R65Cx2.vhd:1275:33  */
  assign n870_o = nextcpucycle == 5'b01100;
  assign n871_o = {n870_o, n864_o, n858_o, n856_o, n854_o, n852_o};
  /* R65Cx2.vhd:1263:33  */
  always @*
    case (n871_o)
      6'b100000: n876_o <= n868_o;
      6'b010000: n876_o <= n862_o;
      6'b001000: n876_o <= 1'b1;
      6'b000100: n876_o <= 1'b1;
      6'b000010: n876_o <= 1'b1;
      6'b000001: n876_o <= n850_o;
    endcase
  /* R65Cx2.vhd:1261:25  */
  assign n878_o = n879_o ? n844_o : s;
  /* R65Cx2.vhd:1261:25  */
  assign n879_o = enable & n876_o;
  /* R65Cx2.vhd:1288:43  */
  assign n881_o = opcinfo[40];
  /* R65Cx2.vhd:1287:25  */
  assign n882_o = n883_o ? aluregisterout : n878_o;
  /* R65Cx2.vhd:1287:25  */
  assign n883_o = updateregisters & n881_o;
  /* R65Cx2.vhd:1253:17  */
  always @(posedge clk)
    n888_q <= n882_o;
  /* R65Cx2.vhd:1305:99  */
  assign n891_o = opcinfo[18];
  /* R65Cx2.vhd:1305:128  */
  assign n892_o = ~irqactive;
  /* R65Cx2.vhd:1305:114  */
  assign n893_o = n891_o & n892_o;
  /* R65Cx2.vhd:1306:148  */
  assign n894_o = myaddrincr[15:8];
  /* R65Cx2.vhd:1308:140  */
  assign n895_o = pc[15:8];
  /* R65Cx2.vhd:1305:89  */
  assign n896_o = n893_o ? n894_o : n895_o;
  /* R65Cx2.vhd:1305:33  */
  assign n898_o = nextcpucycle == 5'b01110;
  /* R65Cx2.vhd:1310:92  */
  assign n899_o = pc[7:0];
  /* R65Cx2.vhd:1310:33  */
  assign n901_o = nextcpucycle == 5'b01111;
  /* R65Cx2.vhd:1311:33  */
  assign n903_o = nextcpucycle == 5'b01010;
  assign n904_o = {n903_o, n901_o, n898_o};
  /* R65Cx2.vhd:1304:33  */
  always @*
    case (n904_o)
      3'b100: n905_o <= di;
      3'b010: n905_o <= n899_o;
      3'b001: n905_o <= n896_o;
    endcase
  /* R65Cx2.vhd:1301:17  */
  assign n909_o = enable ? n905_o : doreg;
  /* R65Cx2.vhd:1301:17  */
  always @(posedge clk)
    n910_q <= n909_o;
  /* R65Cx2.vhd:1331:75  */
  assign n913_o = opcinfo[23];
  /* R65Cx2.vhd:1331:88  */
  assign n914_o = ~n913_o;
  /* R65Cx2.vhd:1331:107  */
  assign n915_o = opcinfo[29];
  /* R65Cx2.vhd:1331:122  */
  assign n916_o = ~n915_o;
  /* R65Cx2.vhd:1331:140  */
  assign n917_o = opcinfo[28];
  /* R65Cx2.vhd:1331:129  */
  assign n918_o = n916_o | n917_o;
  /* R65Cx2.vhd:1331:94  */
  assign n919_o = n914_o & n918_o;
  /* R65Cx2.vhd:1331:65  */
  assign n922_o = n919_o ? 1'b0 : 1'b1;
  /* R65Cx2.vhd:1330:33  */
  assign n924_o = nextcpucycle == 5'b01101;
  /* R65Cx2.vhd:1335:75  */
  assign n925_o = opcinfo[23];
  /* R65Cx2.vhd:1335:88  */
  assign n926_o = ~n925_o;
  /* R65Cx2.vhd:1335:65  */
  assign n929_o = n926_o ? 1'b0 : 1'b1;
  /* R65Cx2.vhd:1334:33  */
  assign n931_o = nextcpucycle == 5'b01110;
  /* R65Cx2.vhd:1334:50  */
  assign n933_o = nextcpucycle == 5'b01111;
  /* R65Cx2.vhd:1334:50  */
  assign n934_o = n931_o | n933_o;
  /* R65Cx2.vhd:1334:64  */
  assign n936_o = nextcpucycle == 5'b10000;
  /* R65Cx2.vhd:1334:64  */
  assign n937_o = n934_o | n936_o;
  /* R65Cx2.vhd:1338:33  */
  assign n939_o = nextcpucycle == 5'b01010;
  /* R65Cx2.vhd:1339:33  */
  assign n941_o = nextcpucycle == 5'b01100;
  assign n942_o = {n941_o, n939_o, n937_o, n924_o};
  /* R65Cx2.vhd:1329:33  */
  always @*
    case (n942_o)
      4'b1000: n946_o <= 1'b0;
      4'b0100: n946_o <= 1'b0;
      4'b0010: n946_o <= n929_o;
      4'b0001: n946_o <= n922_o;
    endcase
  /* R65Cx2.vhd:1326:17  */
  assign n951_o = enable ? n946_o : thewe;
  /* R65Cx2.vhd:1326:17  */
  always @(posedge clk)
    n952_q <= n951_o;
  /* R65Cx2.vhd:1356:33  */
  assign n956_o = thecpucycle == 5'b00000;
  /* R65Cx2.vhd:1357:94  */
  assign n957_o = ~irqactive;
  /* R65Cx2.vhd:1358:123  */
  assign n958_o = opcinfo[33];
  /* R65Cx2.vhd:1358:113  */
  assign n959_o = n958_o ? myaddrincr : myaddr;
  /* R65Cx2.vhd:1357:81  */
  assign n960_o = n957_o ? n959_o : pc;
  /* R65Cx2.vhd:1357:33  */
  assign n962_o = thecpucycle == 5'b00001;
  /* R65Cx2.vhd:1364:91  */
  assign n963_o = opcinfo[32];
  /* R65Cx2.vhd:1364:81  */
  assign n964_o = n963_o ? myaddrincr : pc;
  /* R65Cx2.vhd:1364:33  */
  assign n966_o = thecpucycle == 5'b00010;
  assign n967_o = {n966_o, n962_o, n956_o};
  /* R65Cx2.vhd:1355:33  */
  always @*
    case (n967_o)
      3'b100: n968_o <= n964_o;
      3'b010: n968_o <= n960_o;
      3'b001: n968_o <= myaddr;
    endcase
  /* R65Cx2.vhd:1353:17  */
  assign n972_o = enable ? n968_o : pc;
  /* R65Cx2.vhd:1353:17  */
  always @(posedge clk)
    n973_q <= n972_o;
  /* R65Cx2.vhd:1381:75  */
  assign n975_o = opcinfo[29];
  /* R65Cx2.vhd:1381:106  */
  assign n976_o = opcinfo[28];
  /* R65Cx2.vhd:1381:96  */
  assign n977_o = n975_o | n976_o;
  /* R65Cx2.vhd:1383:102  */
  assign n978_o = opcinfo[32];
  /* R65Cx2.vhd:1385:102  */
  assign n979_o = opcinfo[31];
  /* R65Cx2.vhd:1387:102  */
  assign n980_o = opcinfo[30];
  /* R65Cx2.vhd:1389:102  */
  assign n981_o = opcinfo[33];
  /* R65Cx2.vhd:1389:89  */
  assign n984_o = n981_o ? 4'b0001 : 4'b0000;
  /* R65Cx2.vhd:1387:89  */
  assign n986_o = n980_o ? 4'b1010 : n984_o;
  /* R65Cx2.vhd:1385:89  */
  assign n988_o = n979_o ? 4'b1010 : n986_o;
  /* R65Cx2.vhd:1383:89  */
  assign n990_o = n978_o ? 4'b0001 : n988_o;
  /* R65Cx2.vhd:1381:65  */
  assign n992_o = n977_o ? 4'b1100 : n990_o;
  /* R65Cx2.vhd:1381:17  */
  assign n994_o = thecpucycle == 5'b00001;
  /* R65Cx2.vhd:1394:76  */
  assign n995_o = opcinfo[30];
  /* R65Cx2.vhd:1394:117  */
  assign n996_o = opcinfo[25];
  /* R65Cx2.vhd:1394:105  */
  assign n997_o = n995_o & n996_o;
  /* R65Cx2.vhd:1394:65  */
  assign n1000_o = n997_o ? 4'b1000 : 4'b1001;
  /* R65Cx2.vhd:1394:17  */
  assign n1002_o = thecpucycle == 5'b00010;
  /* R65Cx2.vhd:1399:17  */
  assign n1004_o = thecpucycle == 5'b00011;
  /* R65Cx2.vhd:1400:17  */
  assign n1006_o = thecpucycle == 5'b00100;
  /* R65Cx2.vhd:1401:17  */
  assign n1008_o = thecpucycle == 5'b00101;
  /* R65Cx2.vhd:1402:53  */
  assign n1009_o = t[7];
  /* R65Cx2.vhd:1402:57  */
  assign n1010_o = ~n1009_o;
  /* R65Cx2.vhd:1402:49  */
  assign n1013_o = n1010_o ? 4'b0011 : 4'b0100;
  /* R65Cx2.vhd:1402:17  */
  assign n1015_o = thecpucycle == 5'b00110;
  /* R65Cx2.vhd:1407:17  */
  assign n1017_o = thecpucycle == 5'b00111;
  /* R65Cx2.vhd:1409:99  */
  assign n1018_o = opcinfo[27];
  /* R65Cx2.vhd:1414:103  */
  assign n1019_o = indexout[8];
  /* R65Cx2.vhd:1416:102  */
  assign n1020_o = opcinfo[21];
  /* R65Cx2.vhd:1416:89  */
  assign n1023_o = n1020_o ? 4'b0000 : 4'b0101;
  /* R65Cx2.vhd:1414:89  */
  assign n1025_o = n1019_o ? 4'b0011 : n1023_o;
  /* R65Cx2.vhd:1409:89  */
  assign n1027_o = n1018_o ? 4'b0001 : n1025_o;
  /* R65Cx2.vhd:1408:17  */
  assign n1030_o = thecpucycle == 5'b01000;
  /* R65Cx2.vhd:1420:99  */
  assign n1031_o = opcinfo[21];
  /* R65Cx2.vhd:1420:89  */
  assign n1034_o = n1031_o ? 4'b0000 : 4'b0101;
  /* R65Cx2.vhd:1419:17  */
  assign n1037_o = thecpucycle == 5'b01001;
  /* R65Cx2.vhd:1423:17  */
  assign n1039_o = thecpucycle == 5'b01010;
  /* R65Cx2.vhd:1425:99  */
  assign n1040_o = opcinfo[31];
  /* R65Cx2.vhd:1427:103  */
  assign n1041_o = indexout[8];
  /* R65Cx2.vhd:1427:89  */
  assign n1044_o = n1041_o ? 4'b0011 : 4'b0000;
  /* R65Cx2.vhd:1425:89  */
  assign n1046_o = n1040_o ? 4'b1011 : n1044_o;
  /* R65Cx2.vhd:1424:17  */
  assign n1049_o = thecpucycle == 5'b01011;
  /* R65Cx2.vhd:1430:17  */
  assign n1051_o = thecpucycle == 5'b01100;
  /* R65Cx2.vhd:1431:17  */
  assign n1053_o = thecpucycle == 5'b01101;
  /* R65Cx2.vhd:1432:17  */
  assign n1055_o = thecpucycle == 5'b01110;
  /* R65Cx2.vhd:1434:99  */
  assign n1056_o = opcinfo[28];
  /* R65Cx2.vhd:1434:114  */
  assign n1057_o = ~n1056_o;
  /* R65Cx2.vhd:1434:89  */
  assign n1060_o = n1057_o ? 4'b0101 : 4'b1100;
  /* R65Cx2.vhd:1433:17  */
  assign n1063_o = thecpucycle == 5'b01111;
  /* R65Cx2.vhd:1437:17  */
  assign n1065_o = thecpucycle == 5'b10000;
  /* R65Cx2.vhd:1438:17  */
  assign n1067_o = thecpucycle == 5'b10001;
  assign n1068_o = {n1067_o, n1065_o, n1063_o, n1055_o, n1053_o, n1051_o, n1049_o, n1039_o, n1037_o, n1030_o, n1017_o, n1015_o, n1008_o, n1006_o, n1004_o, n1002_o, n994_o};
  /* R65Cx2.vhd:1380:17  */
  always @*
    case (n1068_o)
      17'b10000000000000000: n1080_o <= 4'b1000;
      17'b01000000000000000: n1080_o <= 4'b0110;
      17'b00100000000000000: n1080_o <= n1060_o;
      17'b00010000000000000: n1080_o <= 4'b1100;
      17'b00001000000000000: n1080_o <= 4'b1100;
      17'b00000100000000000: n1080_o <= 4'b0101;
      17'b00000010000000000: n1080_o <= n1046_o;
      17'b00000001000000000: n1080_o <= 4'b0000;
      17'b00000000100000000: n1080_o <= n1034_o;
      17'b00000000010000000: n1080_o <= n1027_o;
      17'b00000000001000000: n1080_o <= 4'b1011;
      17'b00000000000100000: n1080_o <= n1013_o;
      17'b00000000000010000: n1080_o <= 4'b1101;
      17'b00000000000001000: n1080_o <= 4'b0010;
      17'b00000000000000100: n1080_o <= 4'b1011;
      17'b00000000000000010: n1080_o <= n1000_o;
      17'b00000000000000001: n1080_o <= n992_o;
    endcase
  /* R65Cx2.vhd:1444:26  */
  assign n1082_o = ~reset;
  /* R65Cx2.vhd:1444:17  */
  assign n1084_o = n1082_o ? 4'b0111 : n1080_o;
  /* R65Cx2.vhd:1457:27  */
  assign n1087_o = opcinfo[25];
  /* R65Cx2.vhd:1458:43  */
  assign n1089_o = {1'b0, t};
  /* R65Cx2.vhd:1458:56  */
  assign n1091_o = {1'b0, x};
  /* R65Cx2.vhd:1458:48  */
  assign n1092_o = n1089_o + n1091_o;
  /* R65Cx2.vhd:1459:30  */
  assign n1093_o = opcinfo[24];
  /* R65Cx2.vhd:1460:51  */
  assign n1095_o = {1'b0, t};
  /* R65Cx2.vhd:1460:64  */
  assign n1097_o = {1'b0, y};
  /* R65Cx2.vhd:1460:56  */
  assign n1098_o = n1095_o + n1097_o;
  /* R65Cx2.vhd:1461:30  */
  assign n1099_o = opcinfo[26];
  /* R65Cx2.vhd:1462:43  */
  assign n1101_o = {1'b0, t};
  /* R65Cx2.vhd:1462:64  */
  assign n1102_o = myaddr[7:0];
  /* R65Cx2.vhd:1462:56  */
  assign n1104_o = {1'b0, n1102_o};
  /* R65Cx2.vhd:1462:48  */
  assign n1105_o = n1101_o + n1104_o;
  /* R65Cx2.vhd:1464:42  */
  assign n1107_o = {1'b0, t};
  /* R65Cx2.vhd:1461:17  */
  assign n1108_o = n1099_o ? n1105_o : n1107_o;
  /* R65Cx2.vhd:1459:17  */
  assign n1109_o = n1093_o ? n1098_o : n1108_o;
  /* R65Cx2.vhd:1457:17  */
  assign n1110_o = n1087_o ? n1092_o : n1109_o;
  /* R65Cx2.vhd:1473:33  */
  assign n1115_o = nextaddr == 4'b0001;
  /* R65Cx2.vhd:1474:87  */
  assign n1116_o = myaddrincr[7:0];
  /* R65Cx2.vhd:1474:33  */
  assign n1118_o = nextaddr == 4'b0010;
  /* R65Cx2.vhd:1475:33  */
  assign n1120_o = nextaddr == 4'b0011;
  /* R65Cx2.vhd:1476:33  */
  assign n1122_o = nextaddr == 4'b0100;
  /* R65Cx2.vhd:1477:33  */
  assign n1124_o = nextaddr == 4'b0101;
  /* R65Cx2.vhd:1479:51  */
  assign n1125_o = ~nmireg;
  /* R65Cx2.vhd:1479:41  */
  assign n1128_o = n1125_o ? 16'b1111111111111010 : 16'b1111111111111110;
  /* R65Cx2.vhd:1478:33  */
  assign n1131_o = nextaddr == 4'b0110;
  /* R65Cx2.vhd:1482:33  */
  assign n1133_o = nextaddr == 4'b0111;
  /* R65Cx2.vhd:1483:66  */
  assign n1134_o = {di, t};
  /* R65Cx2.vhd:1483:33  */
  assign n1136_o = nextaddr == 4'b1000;
  /* R65Cx2.vhd:1485:54  */
  assign n1138_o = theopcode == 8'b01111100;
  /* R65Cx2.vhd:1486:63  */
  assign n1139_o = {di, t};
  /* R65Cx2.vhd:1486:76  */
  assign n1141_o = {8'b00000000, x};
  /* R65Cx2.vhd:1486:68  */
  assign n1142_o = n1139_o + n1141_o;
  /* R65Cx2.vhd:1488:72  */
  assign n1143_o = indexout[7:0];
  /* R65Cx2.vhd:1488:62  */
  assign n1144_o = {di, n1143_o};
  /* R65Cx2.vhd:1485:41  */
  assign n1145_o = n1138_o ? n1142_o : n1144_o;
  /* R65Cx2.vhd:1484:33  */
  assign n1147_o = nextaddr == 4'b1001;
  /* R65Cx2.vhd:1490:79  */
  assign n1149_o = {8'b00000000, di};
  /* R65Cx2.vhd:1490:33  */
  assign n1151_o = nextaddr == 4'b1010;
  /* R65Cx2.vhd:1491:90  */
  assign n1152_o = indexout[7:0];
  /* R65Cx2.vhd:1491:80  */
  assign n1154_o = {8'b00000000, n1152_o};
  /* R65Cx2.vhd:1491:33  */
  assign n1156_o = nextaddr == 4'b1011;
  /* R65Cx2.vhd:1492:76  */
  assign n1158_o = {8'b00000001, s};
  /* R65Cx2.vhd:1492:33  */
  assign n1160_o = nextaddr == 4'b1100;
  /* R65Cx2.vhd:1493:88  */
  assign n1161_o = indexout[7:0];
  /* R65Cx2.vhd:1493:33  */
  assign n1163_o = nextaddr == 4'b1101;
  assign n1164_o = {n1163_o, n1160_o, n1156_o, n1151_o, n1147_o, n1136_o, n1133_o, n1131_o, n1124_o, n1122_o, n1120_o, n1118_o, n1115_o};
  assign n1165_o = myaddrincr[7:0];
  assign n1166_o = pc[7:0];
  assign n1167_o = n1128_o[7:0];
  assign n1169_o = n1134_o[7:0];
  assign n1170_o = n1145_o[7:0];
  assign n1171_o = n1149_o[7:0];
  assign n1172_o = n1154_o[7:0];
  assign n1173_o = n1158_o[7:0];
  assign n1174_o = myaddr[7:0];
  /* R65Cx2.vhd:1472:33  */
  always @*
    case (n1164_o)
      13'b1000000000000: n1175_o <= n1161_o;
      13'b0100000000000: n1175_o <= n1173_o;
      13'b0010000000000: n1175_o <= n1172_o;
      13'b0001000000000: n1175_o <= n1171_o;
      13'b0000100000000: n1175_o <= n1170_o;
      13'b0000010000000: n1175_o <= n1169_o;
      13'b0000001000000: n1175_o <= 8'b11111111;
      13'b0000000100000: n1175_o <= n1167_o;
      13'b0000000010000: n1175_o <= n1166_o;
      13'b0000000001000: n1175_o <= n1174_o;
      13'b0000000000100: n1175_o <= n1174_o;
      13'b0000000000010: n1175_o <= n1116_o;
      13'b0000000000001: n1175_o <= n1165_o;
    endcase
  assign n1176_o = myaddrincr[15:8];
  assign n1177_o = pc[15:8];
  assign n1178_o = n1128_o[15:8];
  assign n1180_o = n1134_o[15:8];
  assign n1181_o = n1145_o[15:8];
  assign n1182_o = n1149_o[15:8];
  assign n1183_o = n1154_o[15:8];
  assign n1184_o = n1158_o[15:8];
  assign n1185_o = myaddr[15:8];
  /* R65Cx2.vhd:1472:33  */
  always @*
    case (n1164_o)
      13'b1000000000000: n1186_o <= n1185_o;
      13'b0100000000000: n1186_o <= n1184_o;
      13'b0010000000000: n1186_o <= n1183_o;
      13'b0001000000000: n1186_o <= n1182_o;
      13'b0000100000000: n1186_o <= n1181_o;
      13'b0000010000000: n1186_o <= n1180_o;
      13'b0000001000000: n1186_o <= 8'b11111100;
      13'b0000000100000: n1186_o <= n1178_o;
      13'b0000000010000: n1186_o <= n1177_o;
      13'b0000000001000: n1186_o <= myaddrdecrh;
      13'b0000000000100: n1186_o <= myaddrincrh;
      13'b0000000000010: n1186_o <= n1185_o;
      13'b0000000000001: n1186_o <= n1176_o;
    endcase
  assign n1187_o = {n1186_o, n1175_o};
  /* R65Cx2.vhd:1470:17  */
  assign n1191_o = enable ? n1187_o : myaddr;
  /* R65Cx2.vhd:1470:17  */
  always @(posedge clk)
    n1192_q <= n1191_o;
  /* R65Cx2.vhd:1500:30  */
  assign n1194_o = myaddr + 16'b0000000000000001;
  /* R65Cx2.vhd:1501:30  */
  assign n1195_o = myaddr[15:8];
  /* R65Cx2.vhd:1501:44  */
  assign n1197_o = n1195_o + 8'b00000001;
  /* R65Cx2.vhd:1502:30  */
  assign n1198_o = myaddr[15:8];
  /* R65Cx2.vhd:1502:44  */
  assign n1200_o = n1198_o - 8'b00000001;
  /* R65Cx2.vhd:1518:33  */
  assign n1203_o = thecpucycle == 5'b00000;
  /* R65Cx2.vhd:1518:16  */
  assign n1204_o = n1203_o ? 1'b1 : 1'b0;
  /* R65Cx2.vhd:1522:33  */
  assign n1207_o = {pc, 8'b00000001};
  /* R65Cx2.vhd:1523:23  */
  assign n1208_o = {n1207_o, s};
  /* R65Cx2.vhd:1523:44  */
  assign n1209_o = {n1208_o, n};
  /* R65Cx2.vhd:1524:14  */
  assign n1210_o = {n1209_o, v};
  /* R65Cx2.vhd:1524:18  */
  assign n1211_o = {n1210_o, r};
  /* R65Cx2.vhd:1524:22  */
  assign n1212_o = {n1211_o, b};
  /* R65Cx2.vhd:1524:26  */
  assign n1213_o = {n1212_o, d};
  /* R65Cx2.vhd:1524:30  */
  assign n1214_o = {n1213_o, i};
  /* R65Cx2.vhd:1524:34  */
  assign n1215_o = {n1214_o, z};
  /* R65Cx2.vhd:1524:38  */
  assign n1216_o = {n1215_o, c};
  /* R65Cx2.vhd:1524:42  */
  assign n1217_o = {n1216_o, y};
  /* R65Cx2.vhd:1525:32  */
  assign n1218_o = {n1217_o, x};
  /* R65Cx2.vhd:1526:32  */
  assign n1219_o = {n1218_o, a};
  assign n1223_o = n440_o[43:0];
  assign n1224_o = n440_o[87:44];
  assign n1225_o = n440_o[131:88];
  /* R65Cx2.vhd:31:9  */
  assign n1226_o = n440_o[175:132];
  /* R65Cx2.vhd:29:17  */
  assign n1227_o = n440_o[219:176];
  /* R65Cx2.vhd:28:17  */
  assign n1228_o = n440_o[263:220];
  /* R65Cx2.vhd:27:17  */
  assign n1229_o = n440_o[307:264];
  /* R65Cx2.vhd:26:17  */
  assign n1230_o = n440_o[351:308];
  /* R65Cx2.vhd:25:17  */
  assign n1231_o = n440_o[395:352];
  assign n1232_o = n440_o[439:396];
  assign n1233_o = n440_o[483:440];
  assign n1234_o = n440_o[527:484];
  /* R65Cx2.vhd:1470:17  */
  assign n1235_o = n440_o[571:528];
  assign n1236_o = n440_o[615:572];
  /* R65Cx2.vhd:1468:1  */
  assign n1237_o = n440_o[659:616];
  assign n1238_o = n440_o[703:660];
  /* R65Cx2.vhd:1455:1  */
  assign n1239_o = n440_o[747:704];
  assign n1240_o = n440_o[791:748];
  assign n1241_o = n440_o[835:792];
  assign n1242_o = n440_o[879:836];
  assign n1243_o = n440_o[923:880];
  assign n1244_o = n440_o[967:924];
  assign n1245_o = n440_o[1011:968];
  /* R65Cx2.vhd:1377:1  */
  assign n1246_o = n440_o[1055:1012];
  assign n1247_o = n440_o[1099:1056];
  /* R65Cx2.vhd:1353:17  */
  assign n1248_o = n440_o[1143:1100];
  /* R65Cx2.vhd:1351:1  */
  assign n1249_o = n440_o[1187:1144];
  assign n1250_o = n440_o[1231:1188];
  /* R65Cx2.vhd:1326:17  */
  assign n1251_o = n440_o[1275:1232];
  assign n1252_o = n440_o[1319:1276];
  /* R65Cx2.vhd:1324:1  */
  assign n1253_o = n440_o[1363:1320];
  assign n1254_o = n440_o[1407:1364];
  /* R65Cx2.vhd:1301:17  */
  assign n1255_o = n440_o[1451:1408];
  /* R65Cx2.vhd:1299:1  */
  assign n1256_o = n440_o[1495:1452];
  assign n1257_o = n440_o[1539:1496];
  /* R65Cx2.vhd:1253:17  */
  assign n1258_o = n440_o[1583:1540];
  /* R65Cx2.vhd:1253:17  */
  assign n1259_o = n440_o[1627:1584];
  /* R65Cx2.vhd:1253:17  */
  assign n1260_o = n440_o[1671:1628];
  assign n1261_o = n440_o[1715:1672];
  /* R65Cx2.vhd:1249:9  */
  assign n1262_o = n440_o[1759:1716];
  /* R65Cx2.vhd:1251:26  */
  assign n1263_o = n440_o[1803:1760];
  assign n1264_o = n440_o[1847:1804];
  /* R65Cx2.vhd:1250:26  */
  assign n1265_o = n440_o[1891:1848];
  /* R65Cx2.vhd:1237:17  */
  assign n1266_o = n440_o[1935:1892];
  assign n1267_o = n440_o[1979:1936];
  /* R65Cx2.vhd:1237:17  */
  assign n1268_o = n440_o[2023:1980];
  /* R65Cx2.vhd:1235:9  */
  assign n1269_o = n440_o[2067:2024];
  assign n1270_o = n440_o[2111:2068];
  /* R65Cx2.vhd:1223:17  */
  assign n1271_o = n440_o[2155:2112];
  /* R65Cx2.vhd:1221:9  */
  assign n1272_o = n440_o[2199:2156];
  assign n1273_o = n440_o[2243:2200];
  /* R65Cx2.vhd:1209:9  */
  assign n1274_o = n440_o[2287:2244];
  /* R65Cx2.vhd:1205:9  */
  assign n1275_o = n440_o[2331:2288];
  assign n1276_o = n440_o[2375:2332];
  /* R65Cx2.vhd:1194:9  */
  assign n1277_o = n440_o[2419:2376];
  /* R65Cx2.vhd:1190:9  */
  assign n1278_o = n440_o[2463:2420];
  assign n1279_o = n440_o[2507:2464];
  /* R65Cx2.vhd:1178:17  */
  assign n1280_o = n440_o[2551:2508];
  /* R65Cx2.vhd:1176:9  */
  assign n1281_o = n440_o[2595:2552];
  assign n1282_o = n440_o[2639:2596];
  /* R65Cx2.vhd:1164:17  */
  assign n1283_o = n440_o[2683:2640];
  /* R65Cx2.vhd:1162:9  */
  assign n1284_o = n440_o[2727:2684];
  assign n1285_o = n440_o[2771:2728];
  /* R65Cx2.vhd:1150:17  */
  assign n1286_o = n440_o[2815:2772];
  /* R65Cx2.vhd:1148:9  */
  assign n1287_o = n440_o[2859:2816];
  assign n1288_o = n440_o[2903:2860];
  /* R65Cx2.vhd:1136:17  */
  assign n1289_o = n440_o[2947:2904];
  /* R65Cx2.vhd:1134:9  */
  assign n1290_o = n440_o[2991:2948];
  assign n1291_o = n440_o[3035:2992];
  /* R65Cx2.vhd:1122:17  */
  assign n1292_o = n440_o[3079:3036];
  /* R65Cx2.vhd:1120:9  */
  assign n1293_o = n440_o[3123:3080];
  assign n1294_o = n440_o[3167:3124];
  /* R65Cx2.vhd:1098:17  */
  assign n1295_o = n440_o[3211:3168];
  /* R65Cx2.vhd:1096:1  */
  assign n1296_o = n440_o[3255:3212];
  assign n1297_o = n440_o[3299:3256];
  assign n1298_o = n440_o[3343:3300];
  assign n1299_o = n440_o[3387:3344];
  assign n1300_o = n440_o[3431:3388];
  assign n1301_o = n440_o[3475:3432];
  assign n1302_o = n440_o[3519:3476];
  assign n1303_o = n440_o[3563:3520];
  /* R65Cx2.vhd:982:1  */
  assign n1304_o = n440_o[3607:3564];
  assign n1305_o = n440_o[3651:3608];
  /* R65Cx2.vhd:968:9  */
  assign n1306_o = n440_o[3695:3652];
  assign n1307_o = n440_o[3739:3696];
  assign n1308_o = n440_o[3783:3740];
  /* R65Cx2.vhd:954:9  */
  assign n1309_o = n440_o[3827:3784];
  assign n1310_o = n440_o[3871:3828];
  /* R65Cx2.vhd:937:17  */
  assign n1311_o = n440_o[3915:3872];
  /* R65Cx2.vhd:937:17  */
  assign n1312_o = n440_o[3959:3916];
  assign n1313_o = n440_o[4003:3960];
  /* R65Cx2.vhd:935:1  */
  assign n1314_o = n440_o[4047:4004];
  assign n1315_o = n440_o[4091:4048];
  /* R65Cx2.vhd:926:17  */
  assign n1316_o = n440_o[4135:4092];
  /* R65Cx2.vhd:924:1  */
  assign n1317_o = n440_o[4179:4136];
  /* R65Cx2.vhd:912:40  */
  assign n1318_o = n440_o[4223:4180];
  assign n1319_o = n440_o[4267:4224];
  /* R65Cx2.vhd:898:1  */
  assign n1320_o = n440_o[4311:4268];
  /* R65Cx2.vhd:899:26  */
  assign n1321_o = n440_o[4355:4312];
  /* R65Cx2.vhd:866:17  */
  assign n1322_o = n440_o[4399:4356];
  assign n1323_o = n440_o[4443:4400];
  /* R65Cx2.vhd:866:17  */
  assign n1324_o = n440_o[4487:4444];
  /* R65Cx2.vhd:866:17  */
  assign n1325_o = n440_o[4531:4488];
  /* R65Cx2.vhd:866:17  */
  assign n1326_o = n440_o[4575:4532];
  /* R65Cx2.vhd:866:17  */
  assign n1327_o = n440_o[4619:4576];
  /* R65Cx2.vhd:864:1  */
  assign n1328_o = n440_o[4663:4620];
  assign n1329_o = n440_o[4707:4664];
  assign n1330_o = n440_o[4751:4708];
  assign n1331_o = n440_o[4795:4752];
  assign n1332_o = n440_o[4839:4796];
  assign n1333_o = n440_o[4883:4840];
  assign n1334_o = n440_o[4927:4884];
  assign n1335_o = n440_o[4971:4928];
  assign n1336_o = n440_o[5015:4972];
  /* R65Cx2.vhd:707:1  */
  assign n1337_o = n440_o[5059:5016];
  /* R65Cx2.vhd:716:26  */
  assign n1338_o = n440_o[5103:5060];
  assign n1339_o = n440_o[5147:5104];
  /* R65Cx2.vhd:715:26  */
  assign n1340_o = n440_o[5191:5148];
  assign n1341_o = n440_o[5235:5192];
  /* R65Cx2.vhd:714:26  */
  assign n1342_o = n440_o[5279:5236];
  assign n1343_o = n440_o[5323:5280];
  /* R65Cx2.vhd:713:26  */
  assign n1344_o = n440_o[5367:5324];
  assign n1345_o = n440_o[5411:5368];
  /* R65Cx2.vhd:711:26  */
  assign n1346_o = n440_o[5455:5412];
  assign n1347_o = n440_o[5499:5456];
  /* R65Cx2.vhd:710:26  */
  assign n1348_o = n440_o[5543:5500];
  assign n1349_o = n440_o[5587:5544];
  /* R65Cx2.vhd:709:26  */
  assign n1350_o = n440_o[5631:5588];
  assign n1351_o = n440_o[5675:5632];
  /* R65Cx2.vhd:708:26  */
  assign n1352_o = n440_o[5719:5676];
  assign n1353_o = n440_o[5763:5720];
  assign n1354_o = n440_o[5807:5764];
  assign n1355_o = n440_o[5851:5808];
  /* R65Cx2.vhd:671:1  */
  assign n1356_o = n440_o[5895:5852];
  /* R65Cx2.vhd:672:26  */
  assign n1357_o = n440_o[5939:5896];
  assign n1358_o = n440_o[5983:5940];
  assign n1359_o = n440_o[6027:5984];
  assign n1360_o = n440_o[6071:6028];
  /* R65Cx2.vhd:640:1  */
  assign n1361_o = n440_o[6115:6072];
  /* R65Cx2.vhd:641:26  */
  assign n1362_o = n440_o[6159:6116];
  assign n1363_o = n440_o[6203:6160];
  /* R65Cx2.vhd:638:16  */
  assign n1364_o = n440_o[6247:6204];
  /* R65Cx2.vhd:574:16  */
  assign n1365_o = n440_o[6291:6248];
  /* R65Cx2.vhd:84:16  */
  assign n1366_o = n440_o[6335:6292];
  assign n1367_o = n440_o[6379:6336];
  assign n1368_o = n440_o[6423:6380];
  assign n1369_o = n440_o[6467:6424];
  assign n1370_o = n440_o[6511:6468];
  assign n1371_o = n440_o[6555:6512];
  assign n1372_o = n440_o[6599:6556];
  assign n1373_o = n440_o[6643:6600];
  assign n1374_o = n440_o[6687:6644];
  assign n1375_o = n440_o[6731:6688];
  assign n1376_o = n440_o[6775:6732];
  assign n1377_o = n440_o[6819:6776];
  assign n1378_o = n440_o[6863:6820];
  assign n1379_o = n440_o[6907:6864];
  assign n1380_o = n440_o[6951:6908];
  assign n1381_o = n440_o[6995:6952];
  assign n1382_o = n440_o[7039:6996];
  assign n1383_o = n440_o[7083:7040];
  assign n1384_o = n440_o[7127:7084];
  assign n1385_o = n440_o[7171:7128];
  assign n1386_o = n440_o[7215:7172];
  assign n1387_o = n440_o[7259:7216];
  assign n1388_o = n440_o[7303:7260];
  assign n1389_o = n440_o[7347:7304];
  assign n1390_o = n440_o[7391:7348];
  assign n1391_o = n440_o[7435:7392];
  assign n1392_o = n440_o[7479:7436];
  assign n1393_o = n440_o[7523:7480];
  assign n1394_o = n440_o[7567:7524];
  assign n1395_o = n440_o[7611:7568];
  assign n1396_o = n440_o[7655:7612];
  assign n1397_o = n440_o[7699:7656];
  assign n1398_o = n440_o[7743:7700];
  assign n1399_o = n440_o[7787:7744];
  assign n1400_o = n440_o[7831:7788];
  assign n1401_o = n440_o[7875:7832];
  assign n1402_o = n440_o[7919:7876];
  assign n1403_o = n440_o[7963:7920];
  assign n1404_o = n440_o[8007:7964];
  assign n1405_o = n440_o[8051:8008];
  assign n1406_o = n440_o[8095:8052];
  assign n1407_o = n440_o[8139:8096];
  assign n1408_o = n440_o[8183:8140];
  assign n1409_o = n440_o[8227:8184];
  assign n1410_o = n440_o[8271:8228];
  assign n1411_o = n440_o[8315:8272];
  assign n1412_o = n440_o[8359:8316];
  assign n1413_o = n440_o[8403:8360];
  assign n1414_o = n440_o[8447:8404];
  assign n1415_o = n440_o[8491:8448];
  assign n1416_o = n440_o[8535:8492];
  assign n1417_o = n440_o[8579:8536];
  assign n1418_o = n440_o[8623:8580];
  assign n1419_o = n440_o[8667:8624];
  assign n1420_o = n440_o[8711:8668];
  assign n1421_o = n440_o[8755:8712];
  assign n1422_o = n440_o[8799:8756];
  assign n1423_o = n440_o[8843:8800];
  assign n1424_o = n440_o[8887:8844];
  assign n1425_o = n440_o[8931:8888];
  assign n1426_o = n440_o[8975:8932];
  assign n1427_o = n440_o[9019:8976];
  assign n1428_o = n440_o[9063:9020];
  assign n1429_o = n440_o[9107:9064];
  assign n1430_o = n440_o[9151:9108];
  assign n1431_o = n440_o[9195:9152];
  assign n1432_o = n440_o[9239:9196];
  assign n1433_o = n440_o[9283:9240];
  assign n1434_o = n440_o[9327:9284];
  assign n1435_o = n440_o[9371:9328];
  assign n1436_o = n440_o[9415:9372];
  assign n1437_o = n440_o[9459:9416];
  assign n1438_o = n440_o[9503:9460];
  assign n1439_o = n440_o[9547:9504];
  assign n1440_o = n440_o[9591:9548];
  assign n1441_o = n440_o[9635:9592];
  assign n1442_o = n440_o[9679:9636];
  assign n1443_o = n440_o[9723:9680];
  assign n1444_o = n440_o[9767:9724];
  assign n1445_o = n440_o[9811:9768];
  assign n1446_o = n440_o[9855:9812];
  assign n1447_o = n440_o[9899:9856];
  assign n1448_o = n440_o[9943:9900];
  assign n1449_o = n440_o[9987:9944];
  assign n1450_o = n440_o[10031:9988];
  assign n1451_o = n440_o[10075:10032];
  assign n1452_o = n440_o[10119:10076];
  assign n1453_o = n440_o[10163:10120];
  assign n1454_o = n440_o[10207:10164];
  assign n1455_o = n440_o[10251:10208];
  assign n1456_o = n440_o[10295:10252];
  assign n1457_o = n440_o[10339:10296];
  assign n1458_o = n440_o[10383:10340];
  assign n1459_o = n440_o[10427:10384];
  assign n1460_o = n440_o[10471:10428];
  assign n1461_o = n440_o[10515:10472];
  assign n1462_o = n440_o[10559:10516];
  assign n1463_o = n440_o[10603:10560];
  assign n1464_o = n440_o[10647:10604];
  assign n1465_o = n440_o[10691:10648];
  assign n1466_o = n440_o[10735:10692];
  assign n1467_o = n440_o[10779:10736];
  assign n1468_o = n440_o[10823:10780];
  assign n1469_o = n440_o[10867:10824];
  assign n1470_o = n440_o[10911:10868];
  assign n1471_o = n440_o[10955:10912];
  assign n1472_o = n440_o[10999:10956];
  assign n1473_o = n440_o[11043:11000];
  assign n1474_o = n440_o[11087:11044];
  assign n1475_o = n440_o[11131:11088];
  assign n1476_o = n440_o[11175:11132];
  assign n1477_o = n440_o[11219:11176];
  assign n1478_o = n440_o[11263:11220];
  /* R65Cx2.vhd:912:39  */
  assign n1479_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1479_o)
      2'b00: n1480_o <= n1223_o;
      2'b01: n1480_o <= n1224_o;
      2'b10: n1480_o <= n1225_o;
      2'b11: n1480_o <= n1226_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1481_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1481_o)
      2'b00: n1482_o <= n1227_o;
      2'b01: n1482_o <= n1228_o;
      2'b10: n1482_o <= n1229_o;
      2'b11: n1482_o <= n1230_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1483_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1483_o)
      2'b00: n1484_o <= n1231_o;
      2'b01: n1484_o <= n1232_o;
      2'b10: n1484_o <= n1233_o;
      2'b11: n1484_o <= n1234_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1485_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1485_o)
      2'b00: n1486_o <= n1235_o;
      2'b01: n1486_o <= n1236_o;
      2'b10: n1486_o <= n1237_o;
      2'b11: n1486_o <= n1238_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1487_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1487_o)
      2'b00: n1488_o <= n1239_o;
      2'b01: n1488_o <= n1240_o;
      2'b10: n1488_o <= n1241_o;
      2'b11: n1488_o <= n1242_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1489_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1489_o)
      2'b00: n1490_o <= n1243_o;
      2'b01: n1490_o <= n1244_o;
      2'b10: n1490_o <= n1245_o;
      2'b11: n1490_o <= n1246_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1491_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1491_o)
      2'b00: n1492_o <= n1247_o;
      2'b01: n1492_o <= n1248_o;
      2'b10: n1492_o <= n1249_o;
      2'b11: n1492_o <= n1250_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1493_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1493_o)
      2'b00: n1494_o <= n1251_o;
      2'b01: n1494_o <= n1252_o;
      2'b10: n1494_o <= n1253_o;
      2'b11: n1494_o <= n1254_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1495_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1495_o)
      2'b00: n1496_o <= n1255_o;
      2'b01: n1496_o <= n1256_o;
      2'b10: n1496_o <= n1257_o;
      2'b11: n1496_o <= n1258_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1497_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1497_o)
      2'b00: n1498_o <= n1259_o;
      2'b01: n1498_o <= n1260_o;
      2'b10: n1498_o <= n1261_o;
      2'b11: n1498_o <= n1262_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1499_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1499_o)
      2'b00: n1500_o <= n1263_o;
      2'b01: n1500_o <= n1264_o;
      2'b10: n1500_o <= n1265_o;
      2'b11: n1500_o <= n1266_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1501_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1501_o)
      2'b00: n1502_o <= n1267_o;
      2'b01: n1502_o <= n1268_o;
      2'b10: n1502_o <= n1269_o;
      2'b11: n1502_o <= n1270_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1503_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1503_o)
      2'b00: n1504_o <= n1271_o;
      2'b01: n1504_o <= n1272_o;
      2'b10: n1504_o <= n1273_o;
      2'b11: n1504_o <= n1274_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1505_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1505_o)
      2'b00: n1506_o <= n1275_o;
      2'b01: n1506_o <= n1276_o;
      2'b10: n1506_o <= n1277_o;
      2'b11: n1506_o <= n1278_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1507_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1507_o)
      2'b00: n1508_o <= n1279_o;
      2'b01: n1508_o <= n1280_o;
      2'b10: n1508_o <= n1281_o;
      2'b11: n1508_o <= n1282_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1509_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1509_o)
      2'b00: n1510_o <= n1283_o;
      2'b01: n1510_o <= n1284_o;
      2'b10: n1510_o <= n1285_o;
      2'b11: n1510_o <= n1286_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1511_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1511_o)
      2'b00: n1512_o <= n1287_o;
      2'b01: n1512_o <= n1288_o;
      2'b10: n1512_o <= n1289_o;
      2'b11: n1512_o <= n1290_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1513_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1513_o)
      2'b00: n1514_o <= n1291_o;
      2'b01: n1514_o <= n1292_o;
      2'b10: n1514_o <= n1293_o;
      2'b11: n1514_o <= n1294_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1515_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1515_o)
      2'b00: n1516_o <= n1295_o;
      2'b01: n1516_o <= n1296_o;
      2'b10: n1516_o <= n1297_o;
      2'b11: n1516_o <= n1298_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1517_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1517_o)
      2'b00: n1518_o <= n1299_o;
      2'b01: n1518_o <= n1300_o;
      2'b10: n1518_o <= n1301_o;
      2'b11: n1518_o <= n1302_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1519_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1519_o)
      2'b00: n1520_o <= n1303_o;
      2'b01: n1520_o <= n1304_o;
      2'b10: n1520_o <= n1305_o;
      2'b11: n1520_o <= n1306_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1521_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1521_o)
      2'b00: n1522_o <= n1307_o;
      2'b01: n1522_o <= n1308_o;
      2'b10: n1522_o <= n1309_o;
      2'b11: n1522_o <= n1310_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1523_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1523_o)
      2'b00: n1524_o <= n1311_o;
      2'b01: n1524_o <= n1312_o;
      2'b10: n1524_o <= n1313_o;
      2'b11: n1524_o <= n1314_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1525_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1525_o)
      2'b00: n1526_o <= n1315_o;
      2'b01: n1526_o <= n1316_o;
      2'b10: n1526_o <= n1317_o;
      2'b11: n1526_o <= n1318_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1527_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1527_o)
      2'b00: n1528_o <= n1319_o;
      2'b01: n1528_o <= n1320_o;
      2'b10: n1528_o <= n1321_o;
      2'b11: n1528_o <= n1322_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1529_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1529_o)
      2'b00: n1530_o <= n1323_o;
      2'b01: n1530_o <= n1324_o;
      2'b10: n1530_o <= n1325_o;
      2'b11: n1530_o <= n1326_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1531_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1531_o)
      2'b00: n1532_o <= n1327_o;
      2'b01: n1532_o <= n1328_o;
      2'b10: n1532_o <= n1329_o;
      2'b11: n1532_o <= n1330_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1533_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1533_o)
      2'b00: n1534_o <= n1331_o;
      2'b01: n1534_o <= n1332_o;
      2'b10: n1534_o <= n1333_o;
      2'b11: n1534_o <= n1334_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1535_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1535_o)
      2'b00: n1536_o <= n1335_o;
      2'b01: n1536_o <= n1336_o;
      2'b10: n1536_o <= n1337_o;
      2'b11: n1536_o <= n1338_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1537_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1537_o)
      2'b00: n1538_o <= n1339_o;
      2'b01: n1538_o <= n1340_o;
      2'b10: n1538_o <= n1341_o;
      2'b11: n1538_o <= n1342_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1539_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1539_o)
      2'b00: n1540_o <= n1343_o;
      2'b01: n1540_o <= n1344_o;
      2'b10: n1540_o <= n1345_o;
      2'b11: n1540_o <= n1346_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1541_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1541_o)
      2'b00: n1542_o <= n1347_o;
      2'b01: n1542_o <= n1348_o;
      2'b10: n1542_o <= n1349_o;
      2'b11: n1542_o <= n1350_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1543_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1543_o)
      2'b00: n1544_o <= n1351_o;
      2'b01: n1544_o <= n1352_o;
      2'b10: n1544_o <= n1353_o;
      2'b11: n1544_o <= n1354_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1545_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1545_o)
      2'b00: n1546_o <= n1355_o;
      2'b01: n1546_o <= n1356_o;
      2'b10: n1546_o <= n1357_o;
      2'b11: n1546_o <= n1358_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1547_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1547_o)
      2'b00: n1548_o <= n1359_o;
      2'b01: n1548_o <= n1360_o;
      2'b10: n1548_o <= n1361_o;
      2'b11: n1548_o <= n1362_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1549_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1549_o)
      2'b00: n1550_o <= n1363_o;
      2'b01: n1550_o <= n1364_o;
      2'b10: n1550_o <= n1365_o;
      2'b11: n1550_o <= n1366_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1551_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1551_o)
      2'b00: n1552_o <= n1367_o;
      2'b01: n1552_o <= n1368_o;
      2'b10: n1552_o <= n1369_o;
      2'b11: n1552_o <= n1370_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1553_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1553_o)
      2'b00: n1554_o <= n1371_o;
      2'b01: n1554_o <= n1372_o;
      2'b10: n1554_o <= n1373_o;
      2'b11: n1554_o <= n1374_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1555_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1555_o)
      2'b00: n1556_o <= n1375_o;
      2'b01: n1556_o <= n1376_o;
      2'b10: n1556_o <= n1377_o;
      2'b11: n1556_o <= n1378_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1557_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1557_o)
      2'b00: n1558_o <= n1379_o;
      2'b01: n1558_o <= n1380_o;
      2'b10: n1558_o <= n1381_o;
      2'b11: n1558_o <= n1382_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1559_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1559_o)
      2'b00: n1560_o <= n1383_o;
      2'b01: n1560_o <= n1384_o;
      2'b10: n1560_o <= n1385_o;
      2'b11: n1560_o <= n1386_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1561_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1561_o)
      2'b00: n1562_o <= n1387_o;
      2'b01: n1562_o <= n1388_o;
      2'b10: n1562_o <= n1389_o;
      2'b11: n1562_o <= n1390_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1563_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1563_o)
      2'b00: n1564_o <= n1391_o;
      2'b01: n1564_o <= n1392_o;
      2'b10: n1564_o <= n1393_o;
      2'b11: n1564_o <= n1394_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1565_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1565_o)
      2'b00: n1566_o <= n1395_o;
      2'b01: n1566_o <= n1396_o;
      2'b10: n1566_o <= n1397_o;
      2'b11: n1566_o <= n1398_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1567_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1567_o)
      2'b00: n1568_o <= n1399_o;
      2'b01: n1568_o <= n1400_o;
      2'b10: n1568_o <= n1401_o;
      2'b11: n1568_o <= n1402_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1569_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1569_o)
      2'b00: n1570_o <= n1403_o;
      2'b01: n1570_o <= n1404_o;
      2'b10: n1570_o <= n1405_o;
      2'b11: n1570_o <= n1406_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1571_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1571_o)
      2'b00: n1572_o <= n1407_o;
      2'b01: n1572_o <= n1408_o;
      2'b10: n1572_o <= n1409_o;
      2'b11: n1572_o <= n1410_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1573_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1573_o)
      2'b00: n1574_o <= n1411_o;
      2'b01: n1574_o <= n1412_o;
      2'b10: n1574_o <= n1413_o;
      2'b11: n1574_o <= n1414_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1575_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1575_o)
      2'b00: n1576_o <= n1415_o;
      2'b01: n1576_o <= n1416_o;
      2'b10: n1576_o <= n1417_o;
      2'b11: n1576_o <= n1418_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1577_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1577_o)
      2'b00: n1578_o <= n1419_o;
      2'b01: n1578_o <= n1420_o;
      2'b10: n1578_o <= n1421_o;
      2'b11: n1578_o <= n1422_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1579_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1579_o)
      2'b00: n1580_o <= n1423_o;
      2'b01: n1580_o <= n1424_o;
      2'b10: n1580_o <= n1425_o;
      2'b11: n1580_o <= n1426_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1581_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1581_o)
      2'b00: n1582_o <= n1427_o;
      2'b01: n1582_o <= n1428_o;
      2'b10: n1582_o <= n1429_o;
      2'b11: n1582_o <= n1430_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1583_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1583_o)
      2'b00: n1584_o <= n1431_o;
      2'b01: n1584_o <= n1432_o;
      2'b10: n1584_o <= n1433_o;
      2'b11: n1584_o <= n1434_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1585_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1585_o)
      2'b00: n1586_o <= n1435_o;
      2'b01: n1586_o <= n1436_o;
      2'b10: n1586_o <= n1437_o;
      2'b11: n1586_o <= n1438_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1587_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1587_o)
      2'b00: n1588_o <= n1439_o;
      2'b01: n1588_o <= n1440_o;
      2'b10: n1588_o <= n1441_o;
      2'b11: n1588_o <= n1442_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1589_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1589_o)
      2'b00: n1590_o <= n1443_o;
      2'b01: n1590_o <= n1444_o;
      2'b10: n1590_o <= n1445_o;
      2'b11: n1590_o <= n1446_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1591_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1591_o)
      2'b00: n1592_o <= n1447_o;
      2'b01: n1592_o <= n1448_o;
      2'b10: n1592_o <= n1449_o;
      2'b11: n1592_o <= n1450_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1593_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1593_o)
      2'b00: n1594_o <= n1451_o;
      2'b01: n1594_o <= n1452_o;
      2'b10: n1594_o <= n1453_o;
      2'b11: n1594_o <= n1454_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1595_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1595_o)
      2'b00: n1596_o <= n1455_o;
      2'b01: n1596_o <= n1456_o;
      2'b10: n1596_o <= n1457_o;
      2'b11: n1596_o <= n1458_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1597_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1597_o)
      2'b00: n1598_o <= n1459_o;
      2'b01: n1598_o <= n1460_o;
      2'b10: n1598_o <= n1461_o;
      2'b11: n1598_o <= n1462_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1599_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1599_o)
      2'b00: n1600_o <= n1463_o;
      2'b01: n1600_o <= n1464_o;
      2'b10: n1600_o <= n1465_o;
      2'b11: n1600_o <= n1466_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1601_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1601_o)
      2'b00: n1602_o <= n1467_o;
      2'b01: n1602_o <= n1468_o;
      2'b10: n1602_o <= n1469_o;
      2'b11: n1602_o <= n1470_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1603_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1603_o)
      2'b00: n1604_o <= n1471_o;
      2'b01: n1604_o <= n1472_o;
      2'b10: n1604_o <= n1473_o;
      2'b11: n1604_o <= n1474_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1605_o = n438_o[1:0];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1605_o)
      2'b00: n1606_o <= n1475_o;
      2'b01: n1606_o <= n1476_o;
      2'b10: n1606_o <= n1477_o;
      2'b11: n1606_o <= n1478_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1607_o = n438_o[3:2];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1607_o)
      2'b00: n1608_o <= n1480_o;
      2'b01: n1608_o <= n1482_o;
      2'b10: n1608_o <= n1484_o;
      2'b11: n1608_o <= n1486_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1609_o = n438_o[3:2];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1609_o)
      2'b00: n1610_o <= n1488_o;
      2'b01: n1610_o <= n1490_o;
      2'b10: n1610_o <= n1492_o;
      2'b11: n1610_o <= n1494_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1611_o = n438_o[3:2];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1611_o)
      2'b00: n1612_o <= n1496_o;
      2'b01: n1612_o <= n1498_o;
      2'b10: n1612_o <= n1500_o;
      2'b11: n1612_o <= n1502_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1613_o = n438_o[3:2];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1613_o)
      2'b00: n1614_o <= n1504_o;
      2'b01: n1614_o <= n1506_o;
      2'b10: n1614_o <= n1508_o;
      2'b11: n1614_o <= n1510_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1615_o = n438_o[3:2];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1615_o)
      2'b00: n1616_o <= n1512_o;
      2'b01: n1616_o <= n1514_o;
      2'b10: n1616_o <= n1516_o;
      2'b11: n1616_o <= n1518_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1617_o = n438_o[3:2];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1617_o)
      2'b00: n1618_o <= n1520_o;
      2'b01: n1618_o <= n1522_o;
      2'b10: n1618_o <= n1524_o;
      2'b11: n1618_o <= n1526_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1619_o = n438_o[3:2];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1619_o)
      2'b00: n1620_o <= n1528_o;
      2'b01: n1620_o <= n1530_o;
      2'b10: n1620_o <= n1532_o;
      2'b11: n1620_o <= n1534_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1621_o = n438_o[3:2];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1621_o)
      2'b00: n1622_o <= n1536_o;
      2'b01: n1622_o <= n1538_o;
      2'b10: n1622_o <= n1540_o;
      2'b11: n1622_o <= n1542_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1623_o = n438_o[3:2];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1623_o)
      2'b00: n1624_o <= n1544_o;
      2'b01: n1624_o <= n1546_o;
      2'b10: n1624_o <= n1548_o;
      2'b11: n1624_o <= n1550_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1625_o = n438_o[3:2];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1625_o)
      2'b00: n1626_o <= n1552_o;
      2'b01: n1626_o <= n1554_o;
      2'b10: n1626_o <= n1556_o;
      2'b11: n1626_o <= n1558_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1627_o = n438_o[3:2];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1627_o)
      2'b00: n1628_o <= n1560_o;
      2'b01: n1628_o <= n1562_o;
      2'b10: n1628_o <= n1564_o;
      2'b11: n1628_o <= n1566_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1629_o = n438_o[3:2];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1629_o)
      2'b00: n1630_o <= n1568_o;
      2'b01: n1630_o <= n1570_o;
      2'b10: n1630_o <= n1572_o;
      2'b11: n1630_o <= n1574_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1631_o = n438_o[3:2];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1631_o)
      2'b00: n1632_o <= n1576_o;
      2'b01: n1632_o <= n1578_o;
      2'b10: n1632_o <= n1580_o;
      2'b11: n1632_o <= n1582_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1633_o = n438_o[3:2];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1633_o)
      2'b00: n1634_o <= n1584_o;
      2'b01: n1634_o <= n1586_o;
      2'b10: n1634_o <= n1588_o;
      2'b11: n1634_o <= n1590_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1635_o = n438_o[3:2];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1635_o)
      2'b00: n1636_o <= n1592_o;
      2'b01: n1636_o <= n1594_o;
      2'b10: n1636_o <= n1596_o;
      2'b11: n1636_o <= n1598_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1637_o = n438_o[3:2];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1637_o)
      2'b00: n1638_o <= n1600_o;
      2'b01: n1638_o <= n1602_o;
      2'b10: n1638_o <= n1604_o;
      2'b11: n1638_o <= n1606_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1639_o = n438_o[5:4];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1639_o)
      2'b00: n1640_o <= n1608_o;
      2'b01: n1640_o <= n1610_o;
      2'b10: n1640_o <= n1612_o;
      2'b11: n1640_o <= n1614_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1641_o = n438_o[5:4];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1641_o)
      2'b00: n1642_o <= n1616_o;
      2'b01: n1642_o <= n1618_o;
      2'b10: n1642_o <= n1620_o;
      2'b11: n1642_o <= n1622_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1643_o = n438_o[5:4];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1643_o)
      2'b00: n1644_o <= n1624_o;
      2'b01: n1644_o <= n1626_o;
      2'b10: n1644_o <= n1628_o;
      2'b11: n1644_o <= n1630_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1645_o = n438_o[5:4];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1645_o)
      2'b00: n1646_o <= n1632_o;
      2'b01: n1646_o <= n1634_o;
      2'b10: n1646_o <= n1636_o;
      2'b11: n1646_o <= n1638_o;
    endcase
  /* R65Cx2.vhd:912:39  */
  assign n1647_o = n438_o[7:6];
  /* R65Cx2.vhd:912:39  */
  always @*
    case (n1647_o)
      2'b00: n1648_o <= n1640_o;
      2'b01: n1648_o <= n1642_o;
      2'b10: n1648_o <= n1644_o;
      2'b11: n1648_o <= n1646_o;
    endcase
endmodule

